// SAITO Original //////////////////////////////////////////////////////////////////////////////////

module hsd_divider
(
	input [20:0]  INPUT_0,
	input [20:0]  INPUT_1,

	output [30:0] ANSWER
);


wire [29:0] ex_input0;
wire [29:0] ex_input1;
wire [20:0] comp_input0;
wire [20:0] comp_input1;
wire [30:0] tmp_answer;
// for 20bit
wire [20:0] def_20_0;
wire [20:0] def_20_1;
wire [20:0] def_20_2;
wire [20:0] def_20_3;
wire [20:0] def_20_4;
wire [20:0] def_20_5;
wire [20:0] def_20_6;
wire [20:0] def_20_7;
wire [20:0] def_20_8;
wire [20:0] def_20_9;
wire [20:0] def_20_10;
wire [29:0] ans_20;
// for 19bit
wire [19:0] def_19_0;
wire [19:0] def_19_1;
wire [19:0] def_19_2;
wire [19:0] def_19_3;
wire [19:0] def_19_4;
wire [19:0] def_19_5;
wire [19:0] def_19_6;
wire [19:0] def_19_7;
wire [19:0] def_19_8;
wire [19:0] def_19_9;
wire [19:0] def_19_10;
wire [19:0] def_19_11;
wire [29:0] ans_19;
// for 18bit
wire [18:0] def_18_0;
wire [18:0] def_18_1;
wire [18:0] def_18_2;
wire [18:0] def_18_3;
wire [18:0] def_18_4;
wire [18:0] def_18_5;
wire [18:0] def_18_6;
wire [18:0] def_18_7;
wire [18:0] def_18_8;
wire [18:0] def_18_9;
wire [18:0] def_18_10;
wire [18:0] def_18_11;
wire [18:0] def_18_12;
wire [29:0] ans_18;
// for 17bit
wire [17:0] def_17_0;
wire [17:0] def_17_1;
wire [17:0] def_17_2;
wire [17:0] def_17_3;
wire [17:0] def_17_4;
wire [17:0] def_17_5;
wire [17:0] def_17_6;
wire [17:0] def_17_7;
wire [17:0] def_17_8;
wire [17:0] def_17_9;
wire [17:0] def_17_10;
wire [17:0] def_17_11;
wire [17:0] def_17_12;
wire [17:0] def_17_13;
wire [29:0] ans_17;
// for 16bit
wire [16:0] def_16_0;
wire [16:0] def_16_1;
wire [16:0] def_16_2;
wire [16:0] def_16_3;
wire [16:0] def_16_4;
wire [16:0] def_16_5;
wire [16:0] def_16_6;
wire [16:0] def_16_7;
wire [16:0] def_16_8;
wire [16:0] def_16_9;
wire [16:0] def_16_10;
wire [16:0] def_16_11;
wire [16:0] def_16_12;
wire [16:0] def_16_13;
wire [16:0] def_16_14;
wire [29:0] ans_16;
// for 15bit
wire [15:0] def_15_0;
wire [15:0] def_15_1;
wire [15:0] def_15_2;
wire [15:0] def_15_3;
wire [15:0] def_15_4;
wire [15:0] def_15_5;
wire [15:0] def_15_6;
wire [15:0] def_15_7;
wire [15:0] def_15_8;
wire [15:0] def_15_9;
wire [15:0] def_15_10;
wire [15:0] def_15_11;
wire [15:0] def_15_12;
wire [15:0] def_15_13;
wire [15:0] def_15_14;
wire [15:0] def_15_15;
wire [29:0] ans_15;
// for 14bit
wire [14:0] def_14_0;
wire [14:0] def_14_1;
wire [14:0] def_14_2;
wire [14:0] def_14_3;
wire [14:0] def_14_4;
wire [14:0] def_14_5;
wire [14:0] def_14_6;
wire [14:0] def_14_7;
wire [14:0] def_14_8;
wire [14:0] def_14_9;
wire [14:0] def_14_10;
wire [14:0] def_14_11;
wire [14:0] def_14_12;
wire [14:0] def_14_13;
wire [14:0] def_14_14;
wire [14:0] def_14_15;
wire [14:0] def_14_16;
wire [29:0] ans_14;
// for 13bit
wire [13:0] def_13_0;
wire [13:0] def_13_1;
wire [13:0] def_13_2;
wire [13:0] def_13_3;
wire [13:0] def_13_4;
wire [13:0] def_13_5;
wire [13:0] def_13_6;
wire [13:0] def_13_7;
wire [13:0] def_13_8;
wire [13:0] def_13_9;
wire [13:0] def_13_10;
wire [13:0] def_13_11;
wire [13:0] def_13_12;
wire [13:0] def_13_13;
wire [13:0] def_13_14;
wire [13:0] def_13_15;
wire [13:0] def_13_16;
wire [13:0] def_13_17;
wire [29:0] ans_13;
// for 12bit
wire [12:0] def_12_0;
wire [12:0] def_12_1;
wire [12:0] def_12_2;
wire [12:0] def_12_3;
wire [12:0] def_12_4;
wire [12:0] def_12_5;
wire [12:0] def_12_6;
wire [12:0] def_12_7;
wire [12:0] def_12_8;
wire [12:0] def_12_9;
wire [12:0] def_12_10;
wire [12:0] def_12_11;
wire [12:0] def_12_12;
wire [12:0] def_12_13;
wire [12:0] def_12_14;
wire [12:0] def_12_15;
wire [12:0] def_12_16;
wire [12:0] def_12_17;
wire [12:0] def_12_18;
wire [29:0] ans_12;
// for 11bit
wire [11:0] def_11_0;
wire [11:0] def_11_1;
wire [11:0] def_11_2;
wire [11:0] def_11_3;
wire [11:0] def_11_4;
wire [11:0] def_11_5;
wire [11:0] def_11_6;
wire [11:0] def_11_7;
wire [11:0] def_11_8;
wire [11:0] def_11_9;
wire [11:0] def_11_10;
wire [11:0] def_11_11;
wire [11:0] def_11_12;
wire [11:0] def_11_13;
wire [11:0] def_11_14;
wire [11:0] def_11_15;
wire [11:0] def_11_16;
wire [11:0] def_11_17;
wire [11:0] def_11_18;
wire [11:0] def_11_19;
wire [29:0] ans_11;
// for 10bit
wire [10:0] def_10_0;
wire [10:0] def_10_1;
wire [10:0] def_10_2;
wire [10:0] def_10_3;
wire [10:0] def_10_4;
wire [10:0] def_10_5;
wire [10:0] def_10_6;
wire [10:0] def_10_7;
wire [10:0] def_10_8;
wire [10:0] def_10_9;
wire [10:0] def_10_10;
wire [10:0] def_10_11;
wire [10:0] def_10_12;
wire [10:0] def_10_13;
wire [10:0] def_10_14;
wire [10:0] def_10_15;
wire [10:0] def_10_16;
wire [10:0] def_10_17;
wire [10:0] def_10_18;
wire [10:0] def_10_19;
wire [10:0] def_10_20;
wire [29:0] ans_10;
// for 9bit
wire [ 9:0] def_9_0;
wire [ 9:0] def_9_1;
wire [ 9:0] def_9_2;
wire [ 9:0] def_9_3;
wire [ 9:0] def_9_4;
wire [ 9:0] def_9_5;
wire [ 9:0] def_9_6;
wire [ 9:0] def_9_7;
wire [ 9:0] def_9_8;
wire [ 9:0] def_9_9;
wire [ 9:0] def_9_10;
wire [ 9:0] def_9_11;
wire [ 9:0] def_9_12;
wire [ 9:0] def_9_13;
wire [ 9:0] def_9_14;
wire [ 9:0] def_9_15;
wire [ 9:0] def_9_16;
wire [ 9:0] def_9_17;
wire [ 9:0] def_9_18;
wire [ 9:0] def_9_19;
wire [ 9:0] def_9_20;
wire [ 9:0] def_9_21;
wire [29:0] ans_9;
// for 8bit
wire [ 8:0] def_8_0;
wire [ 8:0] def_8_1;
wire [ 8:0] def_8_2;
wire [ 8:0] def_8_3;
wire [ 8:0] def_8_4;
wire [ 8:0] def_8_5;
wire [ 8:0] def_8_6;
wire [ 8:0] def_8_7;
wire [ 8:0] def_8_8;
wire [ 8:0] def_8_9;
wire [ 8:0] def_8_10;
wire [ 8:0] def_8_11;
wire [ 8:0] def_8_12;
wire [ 8:0] def_8_13;
wire [ 8:0] def_8_14;
wire [ 8:0] def_8_15;
wire [ 8:0] def_8_16;
wire [ 8:0] def_8_17;
wire [ 8:0] def_8_18;
wire [ 8:0] def_8_19;
wire [ 8:0] def_8_20;
wire [ 8:0] def_8_21;
wire [ 8:0] def_8_22;
wire [29:0] ans_8;
// for 7bit
wire [ 7:0] def_7_0;
wire [ 7:0] def_7_1;
wire [ 7:0] def_7_2;
wire [ 7:0] def_7_3;
wire [ 7:0] def_7_4;
wire [ 7:0] def_7_5;
wire [ 7:0] def_7_6;
wire [ 7:0] def_7_7;
wire [ 7:0] def_7_8;
wire [ 7:0] def_7_9;
wire [ 7:0] def_7_10;
wire [ 7:0] def_7_11;
wire [ 7:0] def_7_12;
wire [ 7:0] def_7_13;
wire [ 7:0] def_7_14;
wire [ 7:0] def_7_15;
wire [ 7:0] def_7_16;
wire [ 7:0] def_7_17;
wire [ 7:0] def_7_18;
wire [ 7:0] def_7_19;
wire [ 7:0] def_7_20;
wire [ 7:0] def_7_21;
wire [ 7:0] def_7_22;
wire [ 7:0] def_7_23;
wire [29:0] ans_7;
// for 6bit
wire [ 6:0] def_6_0;
wire [ 6:0] def_6_1;
wire [ 6:0] def_6_2;
wire [ 6:0] def_6_3;
wire [ 6:0] def_6_4;
wire [ 6:0] def_6_5;
wire [ 6:0] def_6_6;
wire [ 6:0] def_6_7;
wire [ 6:0] def_6_8;
wire [ 6:0] def_6_9;
wire [ 6:0] def_6_10;
wire [ 6:0] def_6_11;
wire [ 6:0] def_6_12;
wire [ 6:0] def_6_13;
wire [ 6:0] def_6_14;
wire [ 6:0] def_6_15;
wire [ 6:0] def_6_16;
wire [ 6:0] def_6_17;
wire [ 6:0] def_6_18;
wire [ 6:0] def_6_19;
wire [ 6:0] def_6_20;
wire [ 6:0] def_6_21;
wire [ 6:0] def_6_22;
wire [ 6:0] def_6_23;
wire [ 6:0] def_6_24;
wire [29:0] ans_6;
// for 5bit
wire [ 5:0] def_5_0;
wire [ 5:0] def_5_1;
wire [ 5:0] def_5_2;
wire [ 5:0] def_5_3;
wire [ 5:0] def_5_4;
wire [ 5:0] def_5_5;
wire [ 5:0] def_5_6;
wire [ 5:0] def_5_7;
wire [ 5:0] def_5_8;
wire [ 5:0] def_5_9;
wire [ 5:0] def_5_10;
wire [ 5:0] def_5_11;
wire [ 5:0] def_5_12;
wire [ 5:0] def_5_13;
wire [ 5:0] def_5_14;
wire [ 5:0] def_5_15;
wire [ 5:0] def_5_16;
wire [ 5:0] def_5_17;
wire [ 5:0] def_5_18;
wire [ 5:0] def_5_19;
wire [ 5:0] def_5_20;
wire [ 5:0] def_5_21;
wire [ 5:0] def_5_22;
wire [ 5:0] def_5_23;
wire [ 5:0] def_5_24;
wire [ 5:0] def_5_25;
wire [29:0] ans_5;
// for 4bit
wire [ 4:0] def_4_0;
wire [ 4:0] def_4_1;
wire [ 4:0] def_4_2;
wire [ 4:0] def_4_3;
wire [ 4:0] def_4_4;
wire [ 4:0] def_4_5;
wire [ 4:0] def_4_6;
wire [ 4:0] def_4_7;
wire [ 4:0] def_4_8;
wire [ 4:0] def_4_9;
wire [ 4:0] def_4_10;
wire [ 4:0] def_4_11;
wire [ 4:0] def_4_12;
wire [ 4:0] def_4_13;
wire [ 4:0] def_4_14;
wire [ 4:0] def_4_15;
wire [ 4:0] def_4_16;
wire [ 4:0] def_4_17;
wire [ 4:0] def_4_18;
wire [ 4:0] def_4_19;
wire [ 4:0] def_4_20;
wire [ 4:0] def_4_21;
wire [ 4:0] def_4_22;
wire [ 4:0] def_4_23;
wire [ 4:0] def_4_24;
wire [ 4:0] def_4_25;
wire [ 4:0] def_4_26;
wire [29:0] ans_4;
// for 3bit
wire [ 3:0] def_3_0;
wire [ 3:0] def_3_1;
wire [ 3:0] def_3_2;
wire [ 3:0] def_3_3;
wire [ 3:0] def_3_4;
wire [ 3:0] def_3_5;
wire [ 3:0] def_3_6;
wire [ 3:0] def_3_7;
wire [ 3:0] def_3_8;
wire [ 3:0] def_3_9;
wire [ 3:0] def_3_10;
wire [ 3:0] def_3_11;
wire [ 3:0] def_3_12;
wire [ 3:0] def_3_13;
wire [ 3:0] def_3_14;
wire [ 3:0] def_3_15;
wire [ 3:0] def_3_16;
wire [ 3:0] def_3_17;
wire [ 3:0] def_3_18;
wire [ 3:0] def_3_19;
wire [ 3:0] def_3_20;
wire [ 3:0] def_3_21;
wire [ 3:0] def_3_22;
wire [ 3:0] def_3_23;
wire [ 3:0] def_3_24;
wire [ 3:0] def_3_25;
wire [ 3:0] def_3_26;
wire [ 3:0] def_3_27;
wire [29:0] ans_3;
// for 2bit
wire [ 2:0] def_2_0;
wire [ 2:0] def_2_1;
wire [ 2:0] def_2_2;
wire [ 2:0] def_2_3;
wire [ 2:0] def_2_4;
wire [ 2:0] def_2_5;
wire [ 2:0] def_2_6;
wire [ 2:0] def_2_7;
wire [ 2:0] def_2_8;
wire [ 2:0] def_2_9;
wire [ 2:0] def_2_10;
wire [ 2:0] def_2_11;
wire [ 2:0] def_2_12;
wire [ 2:0] def_2_13;
wire [ 2:0] def_2_14;
wire [ 2:0] def_2_15;
wire [ 2:0] def_2_16;
wire [ 2:0] def_2_17;
wire [ 2:0] def_2_18;
wire [ 2:0] def_2_19;
wire [ 2:0] def_2_20;
wire [ 2:0] def_2_21;
wire [ 2:0] def_2_22;
wire [ 2:0] def_2_23;
wire [ 2:0] def_2_24;
wire [ 2:0] def_2_25;
wire [ 2:0] def_2_26;
wire [ 2:0] def_2_27;
wire [ 2:0] def_2_28;
wire [29:0] ans_2;
// for 1bit
wire [ 1:0] def_1_0;
wire [ 1:0] def_1_1;
wire [ 1:0] def_1_2;
wire [ 1:0] def_1_3;
wire [ 1:0] def_1_4;
wire [ 1:0] def_1_5;
wire [ 1:0] def_1_6;
wire [ 1:0] def_1_7;
wire [ 1:0] def_1_8;
wire [ 1:0] def_1_9;
wire [ 1:0] def_1_10;
wire [ 1:0] def_1_11;
wire [ 1:0] def_1_12;
wire [ 1:0] def_1_13;
wire [ 1:0] def_1_14;
wire [ 1:0] def_1_15;
wire [ 1:0] def_1_16;
wire [ 1:0] def_1_17;
wire [ 1:0] def_1_18;
wire [ 1:0] def_1_19;
wire [ 1:0] def_1_20;
wire [ 1:0] def_1_21;
wire [ 1:0] def_1_22;
wire [ 1:0] def_1_23;
wire [ 1:0] def_1_24;
wire [ 1:0] def_1_25;
wire [ 1:0] def_1_26;
wire [ 1:0] def_1_27;
wire [ 1:0] def_1_28;
wire [ 1:0] def_1_29;
wire [29:0] ans_1;
wire plus;




assign comp_input0 = (~INPUT_0)+1'd1;
assign comp_input1 = (~INPUT_1)+1'd1;
assign ex_input0 = (INPUT_0 << 4'd10)&{5'd30{~INPUT_0[20]}} | (comp_input0<<4'd10)&{5'd30{INPUT_0[20]}};
assign ex_input1 = (INPUT_1 & {5'd30{~INPUT_1[20]}}) | ((comp_input1<<4'd10)&{5'd30{INPUT_1[20]}});

assign plus = ~(INPUT_0[20]^INPUT_1[20]);

// 20bit /////////////////////////////////////////////////////////////////////////////
assign jud_20_0 = ex_input0[29:10] >= ex_input1[19:0];
assign jud_20_1 = ((def_20_0<<1'd1) | ex_input0[9]) >= ex_input1[19:0];
assign jud_20_2 = ((def_20_1<<1'd1) | ex_input0[8]) >= ex_input1[19:0];
assign jud_20_3 = ((def_20_2<<1'd1) | ex_input0[7]) >= ex_input1[19:0];
assign jud_20_4 = ((def_20_3<<1'd1) | ex_input0[6]) >= ex_input1[19:0];
assign jud_20_5 = ((def_20_4<<1'd1) | ex_input0[5]) >= ex_input1[19:0];
assign jud_20_6 = ((def_20_5<<1'd1) | ex_input0[4]) >= ex_input1[19:0];
assign jud_20_7 = ((def_20_6<<1'd1) | ex_input0[3]) >= ex_input1[19:0];
assign jud_20_8 = ((def_20_7<<1'd1) | ex_input0[2]) >= ex_input1[19:0];
assign jud_20_9 = ((def_20_8<<1'd1) | ex_input0[1]) >= ex_input1[19:0];
assign jud_20_10 = ((def_20_9<<1'd1) | ex_input0[0]) >= ex_input1[19:0];

assign def_20_0 = ex_input0[29:10] - (ex_input1[19:0] & {5'd20{jud_20_0}});
assign def_20_1 = ((def_20_0<<1'd1) | ex_input0[9]) - (ex_input1[19:0] & {5'd20{jud_20_1}});
assign def_20_2 = ((def_20_1<<1'd1) | ex_input0[8]) - (ex_input1[19:0] & {5'd20{jud_20_2}});
assign def_20_3 = ((def_20_2<<1'd1) | ex_input0[7]) - (ex_input1[19:0] & {5'd20{jud_20_3}});
assign def_20_4 = ((def_20_3<<1'd1) | ex_input0[6]) - (ex_input1[19:0] & {5'd20{jud_20_4}});
assign def_20_5 = ((def_20_4<<1'd1) | ex_input0[5]) - (ex_input1[19:0] & {5'd20{jud_20_5}});
assign def_20_6 = ((def_20_5<<1'd1) | ex_input0[4]) - (ex_input1[19:0] & {5'd20{jud_20_6}});
assign def_20_7 = ((def_20_6<<1'd1) | ex_input0[3]) - (ex_input1[19:0] & {5'd20{jud_20_7}});
assign def_20_8 = ((def_20_7<<1'd1) | ex_input0[2]) - (ex_input1[19:0] & {5'd20{jud_20_8}});
assign def_20_9 = ((def_20_8<<1'd1) | ex_input0[1]) - (ex_input1[19:0] & {5'd20{jud_20_9}});
assign def_20_10 = ((def_20_9<<1'd1) | ex_input0[0]) - (ex_input1[19:0] & {5'd20{jud_20_10}});

assign ans_20[29] = 1'd0;
assign ans_20[28] = 1'd0;
assign ans_20[27] = 1'd0;
assign ans_20[26] = 1'd0;
assign ans_20[25] = 1'd0;
assign ans_20[24] = 1'd0;
assign ans_20[23] = 1'd0;
assign ans_20[22] = 1'd0;
assign ans_20[21] = 1'd0;
assign ans_20[20] = 1'd0;
assign ans_20[19] = 1'd0;
assign ans_20[18] = 1'd0;
assign ans_20[17] = 1'd0;
assign ans_20[16] = 1'd0;
assign ans_20[15] = 1'd0;
assign ans_20[14] = 1'd0;
assign ans_20[13] = 1'd0;
assign ans_20[12] = 1'd0;
assign ans_20[11] = 1'd0;
assign ans_20[10] = jud_20_0;
assign ans_20[9] = jud_20_1;
assign ans_20[8] = jud_20_2;
assign ans_20[7] = jud_20_3;
assign ans_20[6] = jud_20_4;
assign ans_20[5] = jud_20_5;
assign ans_20[4] = jud_20_6;
assign ans_20[3] = jud_20_7;
assign ans_20[2] = jud_20_8;
assign ans_20[1] = jud_20_9;
assign ans_20[0] = jud_20_10;

// 19bit /////////////////////////////////////////////////////////////////////////////
assign jud_19_0 = ex_input0[29:11] >= ex_input1[18:0];
assign jud_19_1 = ((def_19_0<<1'd1) | ex_input0[10]) >= ex_input1[18:0];
assign jud_19_2 = ((def_19_1<<1'd1) | ex_input0[9]) >= ex_input1[18:0];
assign jud_19_3 = ((def_19_2<<1'd1) | ex_input0[8]) >= ex_input1[18:0];
assign jud_19_4 = ((def_19_3<<1'd1) | ex_input0[7]) >= ex_input1[18:0];
assign jud_19_5 = ((def_19_4<<1'd1) | ex_input0[6]) >= ex_input1[18:0];
assign jud_19_6 = ((def_19_5<<1'd1) | ex_input0[5]) >= ex_input1[18:0];
assign jud_19_7 = ((def_19_6<<1'd1) | ex_input0[4]) >= ex_input1[18:0];
assign jud_19_8 = ((def_19_7<<1'd1) | ex_input0[3]) >= ex_input1[18:0];
assign jud_19_9 = ((def_19_8<<1'd1) | ex_input0[2]) >= ex_input1[18:0];
assign jud_19_10 = ((def_19_9<<1'd1) | ex_input0[1]) >= ex_input1[18:0];
assign jud_19_11 = ((def_19_10<<1'd1) | ex_input0[0]) >= ex_input1[18:0];

assign def_19_0 = ex_input0[29:11] - (ex_input1[18:0] & {5'd19{jud_19_0}});
assign def_19_1 = ((def_19_0<<1'd1) | ex_input0[10]) - (ex_input1[18:0] & {5'd19{jud_19_1}});
assign def_19_2 = ((def_19_1<<1'd1) | ex_input0[9]) - (ex_input1[18:0] & {5'd19{jud_19_2}});
assign def_19_3 = ((def_19_2<<1'd1) | ex_input0[8]) - (ex_input1[18:0] & {5'd19{jud_19_3}});
assign def_19_4 = ((def_19_3<<1'd1) | ex_input0[7]) - (ex_input1[18:0] & {5'd19{jud_19_4}});
assign def_19_5 = ((def_19_4<<1'd1) | ex_input0[6]) - (ex_input1[18:0] & {5'd19{jud_19_5}});
assign def_19_6 = ((def_19_5<<1'd1) | ex_input0[5]) - (ex_input1[18:0] & {5'd19{jud_19_6}});
assign def_19_7 = ((def_19_6<<1'd1) | ex_input0[4]) - (ex_input1[18:0] & {5'd19{jud_19_7}});
assign def_19_8 = ((def_19_7<<1'd1) | ex_input0[3]) - (ex_input1[18:0] & {5'd19{jud_19_8}});
assign def_19_9 = ((def_19_8<<1'd1) | ex_input0[2]) - (ex_input1[18:0] & {5'd19{jud_19_9}});
assign def_19_10 = ((def_19_9<<1'd1) | ex_input0[1]) - (ex_input1[18:0] & {5'd19{jud_19_10}});
assign def_19_11 = ((def_19_10<<1'd1) | ex_input0[0]) - (ex_input1[18:0] & {5'd19{jud_19_11}});

assign ans_19[29] = 1'd0;
assign ans_19[28] = 1'd0;
assign ans_19[27] = 1'd0;
assign ans_19[26] = 1'd0;
assign ans_19[25] = 1'd0;
assign ans_19[24] = 1'd0;
assign ans_19[23] = 1'd0;
assign ans_19[22] = 1'd0;
assign ans_19[21] = 1'd0;
assign ans_19[20] = 1'd0;
assign ans_19[19] = 1'd0;
assign ans_19[18] = 1'd0;
assign ans_19[17] = 1'd0;
assign ans_19[16] = 1'd0;
assign ans_19[15] = 1'd0;
assign ans_19[14] = 1'd0;
assign ans_19[13] = 1'd0;
assign ans_19[12] = 1'd0;
assign ans_19[11] = jud_19_0;
assign ans_19[10] = jud_19_1;
assign ans_19[9] = jud_19_2;
assign ans_19[8] = jud_19_3;
assign ans_19[7] = jud_19_4;
assign ans_19[6] = jud_19_5;
assign ans_19[5] = jud_19_6;
assign ans_19[4] = jud_19_7;
assign ans_19[3] = jud_19_8;
assign ans_19[2] = jud_19_9;
assign ans_19[1] = jud_19_10;
assign ans_19[0] = jud_19_11;

// 18bit /////////////////////////////////////////////////////////////////////////////
assign jud_18_0 = ex_input0[29:12] >= ex_input1[17:0];
assign jud_18_1 = ((def_18_0<<1'd1) | ex_input0[11]) >= ex_input1[17:0];
assign jud_18_2 = ((def_18_1<<1'd1) | ex_input0[10]) >= ex_input1[17:0];
assign jud_18_3 = ((def_18_2<<1'd1) | ex_input0[9]) >= ex_input1[17:0];
assign jud_18_4 = ((def_18_3<<1'd1) | ex_input0[8]) >= ex_input1[17:0];
assign jud_18_5 = ((def_18_4<<1'd1) | ex_input0[7]) >= ex_input1[17:0];
assign jud_18_6 = ((def_18_5<<1'd1) | ex_input0[6]) >= ex_input1[17:0];
assign jud_18_7 = ((def_18_6<<1'd1) | ex_input0[5]) >= ex_input1[17:0];
assign jud_18_8 = ((def_18_7<<1'd1) | ex_input0[4]) >= ex_input1[17:0];
assign jud_18_9 = ((def_18_8<<1'd1) | ex_input0[3]) >= ex_input1[17:0];
assign jud_18_10 = ((def_18_9<<1'd1) | ex_input0[2]) >= ex_input1[17:0];
assign jud_18_11 = ((def_18_10<<1'd1) | ex_input0[1]) >= ex_input1[17:0];
assign jud_18_12 = ((def_18_11<<1'd1) | ex_input0[0]) >= ex_input1[17:0];

assign def_18_0 = ex_input0[29:12] - (ex_input1[17:0] & {5'd18{jud_18_0}});
assign def_18_1 = ((def_18_0<<1'd1) | ex_input0[11]) - (ex_input1[17:0] & {5'd18{jud_18_1}});
assign def_18_2 = ((def_18_1<<1'd1) | ex_input0[10]) - (ex_input1[17:0] & {5'd18{jud_18_2}});
assign def_18_3 = ((def_18_2<<1'd1) | ex_input0[9]) - (ex_input1[17:0] & {5'd18{jud_18_3}});
assign def_18_4 = ((def_18_3<<1'd1) | ex_input0[8]) - (ex_input1[17:0] & {5'd18{jud_18_4}});
assign def_18_5 = ((def_18_4<<1'd1) | ex_input0[7]) - (ex_input1[17:0] & {5'd18{jud_18_5}});
assign def_18_6 = ((def_18_5<<1'd1) | ex_input0[6]) - (ex_input1[17:0] & {5'd18{jud_18_6}});
assign def_18_7 = ((def_18_6<<1'd1) | ex_input0[5]) - (ex_input1[17:0] & {5'd18{jud_18_7}});
assign def_18_8 = ((def_18_7<<1'd1) | ex_input0[4]) - (ex_input1[17:0] & {5'd18{jud_18_8}});
assign def_18_9 = ((def_18_8<<1'd1) | ex_input0[3]) - (ex_input1[17:0] & {5'd18{jud_18_9}});
assign def_18_10 = ((def_18_9<<1'd1) | ex_input0[2]) - (ex_input1[17:0] & {5'd18{jud_18_10}});
assign def_18_11 = ((def_18_10<<1'd1) | ex_input0[1]) - (ex_input1[17:0] & {5'd18{jud_18_11}});
assign def_18_12 = ((def_18_11<<1'd1) | ex_input0[0]) - (ex_input1[17:0] & {5'd18{jud_18_12}});

assign ans_18[29] = 1'd0;
assign ans_18[28] = 1'd0;
assign ans_18[27] = 1'd0;
assign ans_18[26] = 1'd0;
assign ans_18[25] = 1'd0;
assign ans_18[24] = 1'd0;
assign ans_18[23] = 1'd0;
assign ans_18[22] = 1'd0;
assign ans_18[21] = 1'd0;
assign ans_18[20] = 1'd0;
assign ans_18[19] = 1'd0;
assign ans_18[18] = 1'd0;
assign ans_18[17] = 1'd0;
assign ans_18[16] = 1'd0;
assign ans_18[15] = 1'd0;
assign ans_18[14] = 1'd0;
assign ans_18[13] = 1'd0;
assign ans_18[12] = jud_18_0;
assign ans_18[11] = jud_18_1;
assign ans_18[10] = jud_18_2;
assign ans_18[9] = jud_18_3;
assign ans_18[8] = jud_18_4;
assign ans_18[7] = jud_18_5;
assign ans_18[6] = jud_18_6;
assign ans_18[5] = jud_18_7;
assign ans_18[4] = jud_18_8;
assign ans_18[3] = jud_18_9;
assign ans_18[2] = jud_18_10;
assign ans_18[1] = jud_18_11;
assign ans_18[0] = jud_18_12;

// 17bit /////////////////////////////////////////////////////////////////////////////
assign jud_17_0 = ex_input0[29:13] >= ex_input1[16:0];
assign jud_17_1 = ((def_17_0<<1'd1) | ex_input0[12]) >= ex_input1[16:0];
assign jud_17_2 = ((def_17_1<<1'd1) | ex_input0[11]) >= ex_input1[16:0];
assign jud_17_3 = ((def_17_2<<1'd1) | ex_input0[10]) >= ex_input1[16:0];
assign jud_17_4 = ((def_17_3<<1'd1) | ex_input0[9]) >= ex_input1[16:0];
assign jud_17_5 = ((def_17_4<<1'd1) | ex_input0[8]) >= ex_input1[16:0];
assign jud_17_6 = ((def_17_5<<1'd1) | ex_input0[7]) >= ex_input1[16:0];
assign jud_17_7 = ((def_17_6<<1'd1) | ex_input0[6]) >= ex_input1[16:0];
assign jud_17_8 = ((def_17_7<<1'd1) | ex_input0[5]) >= ex_input1[16:0];
assign jud_17_9 = ((def_17_8<<1'd1) | ex_input0[4]) >= ex_input1[16:0];
assign jud_17_10 = ((def_17_9<<1'd1) | ex_input0[3]) >= ex_input1[16:0];
assign jud_17_11 = ((def_17_10<<1'd1) | ex_input0[2]) >= ex_input1[16:0];
assign jud_17_12 = ((def_17_11<<1'd1) | ex_input0[1]) >= ex_input1[16:0];
assign jud_17_13 = ((def_17_12<<1'd1) | ex_input0[0]) >= ex_input1[16:0];

assign def_17_0 = ex_input0[29:13] - (ex_input1[16:0] & {5'd17{jud_17_0}});
assign def_17_1 = ((def_17_0<<1'd1) | ex_input0[12]) - (ex_input1[16:0] & {5'd17{jud_17_1}});
assign def_17_2 = ((def_17_1<<1'd1) | ex_input0[11]) - (ex_input1[16:0] & {5'd17{jud_17_2}});
assign def_17_3 = ((def_17_2<<1'd1) | ex_input0[10]) - (ex_input1[16:0] & {5'd17{jud_17_3}});
assign def_17_4 = ((def_17_3<<1'd1) | ex_input0[9]) - (ex_input1[16:0] & {5'd17{jud_17_4}});
assign def_17_5 = ((def_17_4<<1'd1) | ex_input0[8]) - (ex_input1[16:0] & {5'd17{jud_17_5}});
assign def_17_6 = ((def_17_5<<1'd1) | ex_input0[7]) - (ex_input1[16:0] & {5'd17{jud_17_6}});
assign def_17_7 = ((def_17_6<<1'd1) | ex_input0[6]) - (ex_input1[16:0] & {5'd17{jud_17_7}});
assign def_17_8 = ((def_17_7<<1'd1) | ex_input0[5]) - (ex_input1[16:0] & {5'd17{jud_17_8}});
assign def_17_9 = ((def_17_8<<1'd1) | ex_input0[4]) - (ex_input1[16:0] & {5'd17{jud_17_9}});
assign def_17_10 = ((def_17_9<<1'd1) | ex_input0[3]) - (ex_input1[16:0] & {5'd17{jud_17_10}});
assign def_17_11 = ((def_17_10<<1'd1) | ex_input0[2]) - (ex_input1[16:0] & {5'd17{jud_17_11}});
assign def_17_12 = ((def_17_11<<1'd1) | ex_input0[1]) - (ex_input1[16:0] & {5'd17{jud_17_12}});
assign def_17_13 = ((def_17_12<<1'd1) | ex_input0[0]) - (ex_input1[16:0] & {5'd17{jud_17_13}});

assign ans_17[29] = 1'd0;
assign ans_17[28] = 1'd0;
assign ans_17[27] = 1'd0;
assign ans_17[26] = 1'd0;
assign ans_17[25] = 1'd0;
assign ans_17[24] = 1'd0;
assign ans_17[23] = 1'd0;
assign ans_17[22] = 1'd0;
assign ans_17[21] = 1'd0;
assign ans_17[20] = 1'd0;
assign ans_17[19] = 1'd0;
assign ans_17[18] = 1'd0;
assign ans_17[17] = 1'd0;
assign ans_17[16] = 1'd0;
assign ans_17[15] = 1'd0;
assign ans_17[14] = 1'd0;
assign ans_17[13] = jud_17_0;
assign ans_17[12] = jud_17_1;
assign ans_17[11] = jud_17_2;
assign ans_17[10] = jud_17_3;
assign ans_17[9] = jud_17_4;
assign ans_17[8] = jud_17_5;
assign ans_17[7] = jud_17_6;
assign ans_17[6] = jud_17_7;
assign ans_17[5] = jud_17_8;
assign ans_17[4] = jud_17_9;
assign ans_17[3] = jud_17_10;
assign ans_17[2] = jud_17_11;
assign ans_17[1] = jud_17_12;
assign ans_17[0] = jud_17_13;

// 16bit /////////////////////////////////////////////////////////////////////////////
assign jud_16_0 = ex_input0[29:14] >= ex_input1[15:0];
assign jud_16_1 = ((def_16_0<<1'd1) | ex_input0[13]) >= ex_input1[15:0];
assign jud_16_2 = ((def_16_1<<1'd1) | ex_input0[12]) >= ex_input1[15:0];
assign jud_16_3 = ((def_16_2<<1'd1) | ex_input0[11]) >= ex_input1[15:0];
assign jud_16_4 = ((def_16_3<<1'd1) | ex_input0[10]) >= ex_input1[15:0];
assign jud_16_5 = ((def_16_4<<1'd1) | ex_input0[9]) >= ex_input1[15:0];
assign jud_16_6 = ((def_16_5<<1'd1) | ex_input0[8]) >= ex_input1[15:0];
assign jud_16_7 = ((def_16_6<<1'd1) | ex_input0[7]) >= ex_input1[15:0];
assign jud_16_8 = ((def_16_7<<1'd1) | ex_input0[6]) >= ex_input1[15:0];
assign jud_16_9 = ((def_16_8<<1'd1) | ex_input0[5]) >= ex_input1[15:0];
assign jud_16_10 = ((def_16_9<<1'd1) | ex_input0[4]) >= ex_input1[15:0];
assign jud_16_11 = ((def_16_10<<1'd1) | ex_input0[3]) >= ex_input1[15:0];
assign jud_16_12 = ((def_16_11<<1'd1) | ex_input0[2]) >= ex_input1[15:0];
assign jud_16_13 = ((def_16_12<<1'd1) | ex_input0[1]) >= ex_input1[15:0];
assign jud_16_14 = ((def_16_13<<1'd1) | ex_input0[0]) >= ex_input1[15:0];

assign def_16_0 = ex_input0[29:14] - (ex_input1[15:0] & {5'd16{jud_16_0}});
assign def_16_1 = ((def_16_0<<1'd1) | ex_input0[13]) - (ex_input1[15:0] & {5'd16{jud_16_1}});
assign def_16_2 = ((def_16_1<<1'd1) | ex_input0[12]) - (ex_input1[15:0] & {5'd16{jud_16_2}});
assign def_16_3 = ((def_16_2<<1'd1) | ex_input0[11]) - (ex_input1[15:0] & {5'd16{jud_16_3}});
assign def_16_4 = ((def_16_3<<1'd1) | ex_input0[10]) - (ex_input1[15:0] & {5'd16{jud_16_4}});
assign def_16_5 = ((def_16_4<<1'd1) | ex_input0[9]) - (ex_input1[15:0] & {5'd16{jud_16_5}});
assign def_16_6 = ((def_16_5<<1'd1) | ex_input0[8]) - (ex_input1[15:0] & {5'd16{jud_16_6}});
assign def_16_7 = ((def_16_6<<1'd1) | ex_input0[7]) - (ex_input1[15:0] & {5'd16{jud_16_7}});
assign def_16_8 = ((def_16_7<<1'd1) | ex_input0[6]) - (ex_input1[15:0] & {5'd16{jud_16_8}});
assign def_16_9 = ((def_16_8<<1'd1) | ex_input0[5]) - (ex_input1[15:0] & {5'd16{jud_16_9}});
assign def_16_10 = ((def_16_9<<1'd1) | ex_input0[4]) - (ex_input1[15:0] & {5'd16{jud_16_10}});
assign def_16_11 = ((def_16_10<<1'd1) | ex_input0[3]) - (ex_input1[15:0] & {5'd16{jud_16_11}});
assign def_16_12 = ((def_16_11<<1'd1) | ex_input0[2]) - (ex_input1[15:0] & {5'd16{jud_16_12}});
assign def_16_13 = ((def_16_12<<1'd1) | ex_input0[1]) - (ex_input1[15:0] & {5'd16{jud_16_13}});
assign def_16_14 = ((def_16_13<<1'd1) | ex_input0[0]) - (ex_input1[15:0] & {5'd16{jud_16_14}});

assign ans_16[29] = 1'd0;
assign ans_16[28] = 1'd0;
assign ans_16[27] = 1'd0;
assign ans_16[26] = 1'd0;
assign ans_16[25] = 1'd0;
assign ans_16[24] = 1'd0;
assign ans_16[23] = 1'd0;
assign ans_16[22] = 1'd0;
assign ans_16[21] = 1'd0;
assign ans_16[20] = 1'd0;
assign ans_16[19] = 1'd0;
assign ans_16[18] = 1'd0;
assign ans_16[17] = 1'd0;
assign ans_16[16] = 1'd0;
assign ans_16[15] = 1'd0;
assign ans_16[14] = jud_16_0;
assign ans_16[13] = jud_16_1;
assign ans_16[12] = jud_16_2;
assign ans_16[11] = jud_16_3;
assign ans_16[10] = jud_16_4;
assign ans_16[9] = jud_16_5;
assign ans_16[8] = jud_16_6;
assign ans_16[7] = jud_16_7;
assign ans_16[6] = jud_16_8;
assign ans_16[5] = jud_16_9;
assign ans_16[4] = jud_16_10;
assign ans_16[3] = jud_16_11;
assign ans_16[2] = jud_16_12;
assign ans_16[1] = jud_16_13;
assign ans_16[0] = jud_16_14;

// 15bit /////////////////////////////////////////////////////////////////////////////
assign jud_15_0 = ex_input0[29:15] >= ex_input1[14:0];
assign jud_15_1 = ((def_15_0<<1'd1) | ex_input0[14]) >= ex_input1[14:0];
assign jud_15_2 = ((def_15_1<<1'd1) | ex_input0[13]) >= ex_input1[14:0];
assign jud_15_3 = ((def_15_2<<1'd1) | ex_input0[12]) >= ex_input1[14:0];
assign jud_15_4 = ((def_15_3<<1'd1) | ex_input0[11]) >= ex_input1[14:0];
assign jud_15_5 = ((def_15_4<<1'd1) | ex_input0[10]) >= ex_input1[14:0];
assign jud_15_6 = ((def_15_5<<1'd1) | ex_input0[9]) >= ex_input1[14:0];
assign jud_15_7 = ((def_15_6<<1'd1) | ex_input0[8]) >= ex_input1[14:0];
assign jud_15_8 = ((def_15_7<<1'd1) | ex_input0[7]) >= ex_input1[14:0];
assign jud_15_9 = ((def_15_8<<1'd1) | ex_input0[6]) >= ex_input1[14:0];
assign jud_15_10 = ((def_15_9<<1'd1) | ex_input0[5]) >= ex_input1[14:0];
assign jud_15_11 = ((def_15_10<<1'd1) | ex_input0[4]) >= ex_input1[14:0];
assign jud_15_12 = ((def_15_11<<1'd1) | ex_input0[3]) >= ex_input1[14:0];
assign jud_15_13 = ((def_15_12<<1'd1) | ex_input0[2]) >= ex_input1[14:0];
assign jud_15_14 = ((def_15_13<<1'd1) | ex_input0[1]) >= ex_input1[14:0];
assign jud_15_15 = ((def_15_14<<1'd1) | ex_input0[0]) >= ex_input1[14:0];

assign def_15_0 = ex_input0[29:15] - (ex_input1[14:0] & {5'd15{jud_15_0}});
assign def_15_1 = ((def_15_0<<1'd1) | ex_input0[14]) - (ex_input1[14:0] & {5'd15{jud_15_1}});
assign def_15_2 = ((def_15_1<<1'd1) | ex_input0[13]) - (ex_input1[14:0] & {5'd15{jud_15_2}});
assign def_15_3 = ((def_15_2<<1'd1) | ex_input0[12]) - (ex_input1[14:0] & {5'd15{jud_15_3}});
assign def_15_4 = ((def_15_3<<1'd1) | ex_input0[11]) - (ex_input1[14:0] & {5'd15{jud_15_4}});
assign def_15_5 = ((def_15_4<<1'd1) | ex_input0[10]) - (ex_input1[14:0] & {5'd15{jud_15_5}});
assign def_15_6 = ((def_15_5<<1'd1) | ex_input0[9]) - (ex_input1[14:0] & {5'd15{jud_15_6}});
assign def_15_7 = ((def_15_6<<1'd1) | ex_input0[8]) - (ex_input1[14:0] & {5'd15{jud_15_7}});
assign def_15_8 = ((def_15_7<<1'd1) | ex_input0[7]) - (ex_input1[14:0] & {5'd15{jud_15_8}});
assign def_15_9 = ((def_15_8<<1'd1) | ex_input0[6]) - (ex_input1[14:0] & {5'd15{jud_15_9}});
assign def_15_10 = ((def_15_9<<1'd1) | ex_input0[5]) - (ex_input1[14:0] & {5'd15{jud_15_10}});
assign def_15_11 = ((def_15_10<<1'd1) | ex_input0[4]) - (ex_input1[14:0] & {5'd15{jud_15_11}});
assign def_15_12 = ((def_15_11<<1'd1) | ex_input0[3]) - (ex_input1[14:0] & {5'd15{jud_15_12}});
assign def_15_13 = ((def_15_12<<1'd1) | ex_input0[2]) - (ex_input1[14:0] & {5'd15{jud_15_13}});
assign def_15_14 = ((def_15_13<<1'd1) | ex_input0[1]) - (ex_input1[14:0] & {5'd15{jud_15_14}});
assign def_15_15 = ((def_15_14<<1'd1) | ex_input0[0]) - (ex_input1[14:0] & {5'd15{jud_15_15}});

assign ans_15[29] = 1'd0;
assign ans_15[28] = 1'd0;
assign ans_15[27] = 1'd0;
assign ans_15[26] = 1'd0;
assign ans_15[25] = 1'd0;
assign ans_15[24] = 1'd0;
assign ans_15[23] = 1'd0;
assign ans_15[22] = 1'd0;
assign ans_15[21] = 1'd0;
assign ans_15[20] = 1'd0;
assign ans_15[19] = 1'd0;
assign ans_15[18] = 1'd0;
assign ans_15[17] = 1'd0;
assign ans_15[16] = 1'd0;
assign ans_15[15] = jud_15_0;
assign ans_15[14] = jud_15_1;
assign ans_15[13] = jud_15_2;
assign ans_15[12] = jud_15_3;
assign ans_15[11] = jud_15_4;
assign ans_15[10] = jud_15_5;
assign ans_15[9] = jud_15_6;
assign ans_15[8] = jud_15_7;
assign ans_15[7] = jud_15_8;
assign ans_15[6] = jud_15_9;
assign ans_15[5] = jud_15_10;
assign ans_15[4] = jud_15_11;
assign ans_15[3] = jud_15_12;
assign ans_15[2] = jud_15_13;
assign ans_15[1] = jud_15_14;
assign ans_15[0] = jud_15_15;

// 14bit /////////////////////////////////////////////////////////////////////////////
assign jud_14_0 = ex_input0[29:16] >= ex_input1[13:0];
assign jud_14_1 = ((def_14_0<<1'd1) | ex_input0[15]) >= ex_input1[13:0];
assign jud_14_2 = ((def_14_1<<1'd1) | ex_input0[14]) >= ex_input1[13:0];
assign jud_14_3 = ((def_14_2<<1'd1) | ex_input0[13]) >= ex_input1[13:0];
assign jud_14_4 = ((def_14_3<<1'd1) | ex_input0[12]) >= ex_input1[13:0];
assign jud_14_5 = ((def_14_4<<1'd1) | ex_input0[11]) >= ex_input1[13:0];
assign jud_14_6 = ((def_14_5<<1'd1) | ex_input0[10]) >= ex_input1[13:0];
assign jud_14_7 = ((def_14_6<<1'd1) | ex_input0[9]) >= ex_input1[13:0];
assign jud_14_8 = ((def_14_7<<1'd1) | ex_input0[8]) >= ex_input1[13:0];
assign jud_14_9 = ((def_14_8<<1'd1) | ex_input0[7]) >= ex_input1[13:0];
assign jud_14_10 = ((def_14_9<<1'd1) | ex_input0[6]) >= ex_input1[13:0];
assign jud_14_11 = ((def_14_10<<1'd1) | ex_input0[5]) >= ex_input1[13:0];
assign jud_14_12 = ((def_14_11<<1'd1) | ex_input0[4]) >= ex_input1[13:0];
assign jud_14_13 = ((def_14_12<<1'd1) | ex_input0[3]) >= ex_input1[13:0];
assign jud_14_14 = ((def_14_13<<1'd1) | ex_input0[2]) >= ex_input1[13:0];
assign jud_14_15 = ((def_14_14<<1'd1) | ex_input0[1]) >= ex_input1[13:0];
assign jud_14_16 = ((def_14_15<<1'd1) | ex_input0[0]) >= ex_input1[13:0];

assign def_14_0 = ex_input0[29:16] - (ex_input1[13:0] & {5'd14{jud_14_0}});
assign def_14_1 = ((def_14_0<<1'd1) | ex_input0[15]) - (ex_input1[13:0] & {5'd14{jud_14_1}});
assign def_14_2 = ((def_14_1<<1'd1) | ex_input0[14]) - (ex_input1[13:0] & {5'd14{jud_14_2}});
assign def_14_3 = ((def_14_2<<1'd1) | ex_input0[13]) - (ex_input1[13:0] & {5'd14{jud_14_3}});
assign def_14_4 = ((def_14_3<<1'd1) | ex_input0[12]) - (ex_input1[13:0] & {5'd14{jud_14_4}});
assign def_14_5 = ((def_14_4<<1'd1) | ex_input0[11]) - (ex_input1[13:0] & {5'd14{jud_14_5}});
assign def_14_6 = ((def_14_5<<1'd1) | ex_input0[10]) - (ex_input1[13:0] & {5'd14{jud_14_6}});
assign def_14_7 = ((def_14_6<<1'd1) | ex_input0[9]) - (ex_input1[13:0] & {5'd14{jud_14_7}});
assign def_14_8 = ((def_14_7<<1'd1) | ex_input0[8]) - (ex_input1[13:0] & {5'd14{jud_14_8}});
assign def_14_9 = ((def_14_8<<1'd1) | ex_input0[7]) - (ex_input1[13:0] & {5'd14{jud_14_9}});
assign def_14_10 = ((def_14_9<<1'd1) | ex_input0[6]) - (ex_input1[13:0] & {5'd14{jud_14_10}});
assign def_14_11 = ((def_14_10<<1'd1) | ex_input0[5]) - (ex_input1[13:0] & {5'd14{jud_14_11}});
assign def_14_12 = ((def_14_11<<1'd1) | ex_input0[4]) - (ex_input1[13:0] & {5'd14{jud_14_12}});
assign def_14_13 = ((def_14_12<<1'd1) | ex_input0[3]) - (ex_input1[13:0] & {5'd14{jud_14_13}});
assign def_14_14 = ((def_14_13<<1'd1) | ex_input0[2]) - (ex_input1[13:0] & {5'd14{jud_14_14}});
assign def_14_15 = ((def_14_14<<1'd1) | ex_input0[1]) - (ex_input1[13:0] & {5'd14{jud_14_15}});
assign def_14_16 = ((def_14_15<<1'd1) | ex_input0[0]) - (ex_input1[13:0] & {5'd14{jud_14_16}});

assign ans_14[29] = 1'd0;
assign ans_14[28] = 1'd0;
assign ans_14[27] = 1'd0;
assign ans_14[26] = 1'd0;
assign ans_14[25] = 1'd0;
assign ans_14[24] = 1'd0;
assign ans_14[23] = 1'd0;
assign ans_14[22] = 1'd0;
assign ans_14[21] = 1'd0;
assign ans_14[20] = 1'd0;
assign ans_14[19] = 1'd0;
assign ans_14[18] = 1'd0;
assign ans_14[17] = 1'd0;
assign ans_14[16] = jud_14_0;
assign ans_14[15] = jud_14_1;
assign ans_14[14] = jud_14_2;
assign ans_14[13] = jud_14_3;
assign ans_14[12] = jud_14_4;
assign ans_14[11] = jud_14_5;
assign ans_14[10] = jud_14_6;
assign ans_14[9] = jud_14_7;
assign ans_14[8] = jud_14_8;
assign ans_14[7] = jud_14_9;
assign ans_14[6] = jud_14_10;
assign ans_14[5] = jud_14_11;
assign ans_14[4] = jud_14_12;
assign ans_14[3] = jud_14_13;
assign ans_14[2] = jud_14_14;
assign ans_14[1] = jud_14_15;
assign ans_14[0] = jud_14_16;

// 13bit /////////////////////////////////////////////////////////////////////////////
assign jud_13_0 = ex_input0[29:17] >= ex_input1[12:0];
assign jud_13_1 = ((def_13_0<<1'd1) | ex_input0[16]) >= ex_input1[12:0];
assign jud_13_2 = ((def_13_1<<1'd1) | ex_input0[15]) >= ex_input1[12:0];
assign jud_13_3 = ((def_13_2<<1'd1) | ex_input0[14]) >= ex_input1[12:0];
assign jud_13_4 = ((def_13_3<<1'd1) | ex_input0[13]) >= ex_input1[12:0];
assign jud_13_5 = ((def_13_4<<1'd1) | ex_input0[12]) >= ex_input1[12:0];
assign jud_13_6 = ((def_13_5<<1'd1) | ex_input0[11]) >= ex_input1[12:0];
assign jud_13_7 = ((def_13_6<<1'd1) | ex_input0[10]) >= ex_input1[12:0];
assign jud_13_8 = ((def_13_7<<1'd1) | ex_input0[9]) >= ex_input1[12:0];
assign jud_13_9 = ((def_13_8<<1'd1) | ex_input0[8]) >= ex_input1[12:0];
assign jud_13_10 = ((def_13_9<<1'd1) | ex_input0[7]) >= ex_input1[12:0];
assign jud_13_11 = ((def_13_10<<1'd1) | ex_input0[6]) >= ex_input1[12:0];
assign jud_13_12 = ((def_13_11<<1'd1) | ex_input0[5]) >= ex_input1[12:0];
assign jud_13_13 = ((def_13_12<<1'd1) | ex_input0[4]) >= ex_input1[12:0];
assign jud_13_14 = ((def_13_13<<1'd1) | ex_input0[3]) >= ex_input1[12:0];
assign jud_13_15 = ((def_13_14<<1'd1) | ex_input0[2]) >= ex_input1[12:0];
assign jud_13_16 = ((def_13_15<<1'd1) | ex_input0[1]) >= ex_input1[12:0];
assign jud_13_17 = ((def_13_16<<1'd1) | ex_input0[0]) >= ex_input1[12:0];

assign def_13_0 = ex_input0[29:17] - (ex_input1[12:0] & {5'd13{jud_13_0}});
assign def_13_1 = ((def_13_0<<1'd1) | ex_input0[16]) - (ex_input1[12:0] & {5'd13{jud_13_1}});
assign def_13_2 = ((def_13_1<<1'd1) | ex_input0[15]) - (ex_input1[12:0] & {5'd13{jud_13_2}});
assign def_13_3 = ((def_13_2<<1'd1) | ex_input0[14]) - (ex_input1[12:0] & {5'd13{jud_13_3}});
assign def_13_4 = ((def_13_3<<1'd1) | ex_input0[13]) - (ex_input1[12:0] & {5'd13{jud_13_4}});
assign def_13_5 = ((def_13_4<<1'd1) | ex_input0[12]) - (ex_input1[12:0] & {5'd13{jud_13_5}});
assign def_13_6 = ((def_13_5<<1'd1) | ex_input0[11]) - (ex_input1[12:0] & {5'd13{jud_13_6}});
assign def_13_7 = ((def_13_6<<1'd1) | ex_input0[10]) - (ex_input1[12:0] & {5'd13{jud_13_7}});
assign def_13_8 = ((def_13_7<<1'd1) | ex_input0[9]) - (ex_input1[12:0] & {5'd13{jud_13_8}});
assign def_13_9 = ((def_13_8<<1'd1) | ex_input0[8]) - (ex_input1[12:0] & {5'd13{jud_13_9}});
assign def_13_10 = ((def_13_9<<1'd1) | ex_input0[7]) - (ex_input1[12:0] & {5'd13{jud_13_10}});
assign def_13_11 = ((def_13_10<<1'd1) | ex_input0[6]) - (ex_input1[12:0] & {5'd13{jud_13_11}});
assign def_13_12 = ((def_13_11<<1'd1) | ex_input0[5]) - (ex_input1[12:0] & {5'd13{jud_13_12}});
assign def_13_13 = ((def_13_12<<1'd1) | ex_input0[4]) - (ex_input1[12:0] & {5'd13{jud_13_13}});
assign def_13_14 = ((def_13_13<<1'd1) | ex_input0[3]) - (ex_input1[12:0] & {5'd13{jud_13_14}});
assign def_13_15 = ((def_13_14<<1'd1) | ex_input0[2]) - (ex_input1[12:0] & {5'd13{jud_13_15}});
assign def_13_16 = ((def_13_15<<1'd1) | ex_input0[1]) - (ex_input1[12:0] & {5'd13{jud_13_16}});
assign def_13_17 = ((def_13_16<<1'd1) | ex_input0[0]) - (ex_input1[12:0] & {5'd13{jud_13_17}});

assign ans_13[29] = 1'd0;
assign ans_13[28] = 1'd0;
assign ans_13[27] = 1'd0;
assign ans_13[26] = 1'd0;
assign ans_13[25] = 1'd0;
assign ans_13[24] = 1'd0;
assign ans_13[23] = 1'd0;
assign ans_13[22] = 1'd0;
assign ans_13[21] = 1'd0;
assign ans_13[20] = 1'd0;
assign ans_13[19] = 1'd0;
assign ans_13[18] = 1'd0;
assign ans_13[17] = jud_13_0;
assign ans_13[16] = jud_13_1;
assign ans_13[15] = jud_13_2;
assign ans_13[14] = jud_13_3;
assign ans_13[13] = jud_13_4;
assign ans_13[12] = jud_13_5;
assign ans_13[11] = jud_13_6;
assign ans_13[10] = jud_13_7;
assign ans_13[9] = jud_13_8;
assign ans_13[8] = jud_13_9;
assign ans_13[7] = jud_13_10;
assign ans_13[6] = jud_13_11;
assign ans_13[5] = jud_13_12;
assign ans_13[4] = jud_13_13;
assign ans_13[3] = jud_13_14;
assign ans_13[2] = jud_13_15;
assign ans_13[1] = jud_13_16;
assign ans_13[0] = jud_13_17;

// 12bit /////////////////////////////////////////////////////////////////////////////
assign jud_12_0 = ex_input0[29:18] >= ex_input1[11:0];
assign jud_12_1 = ((def_12_0<<1'd1) | ex_input0[17]) >= ex_input1[11:0];
assign jud_12_2 = ((def_12_1<<1'd1) | ex_input0[16]) >= ex_input1[11:0];
assign jud_12_3 = ((def_12_2<<1'd1) | ex_input0[15]) >= ex_input1[11:0];
assign jud_12_4 = ((def_12_3<<1'd1) | ex_input0[14]) >= ex_input1[11:0];
assign jud_12_5 = ((def_12_4<<1'd1) | ex_input0[13]) >= ex_input1[11:0];
assign jud_12_6 = ((def_12_5<<1'd1) | ex_input0[12]) >= ex_input1[11:0];
assign jud_12_7 = ((def_12_6<<1'd1) | ex_input0[11]) >= ex_input1[11:0];
assign jud_12_8 = ((def_12_7<<1'd1) | ex_input0[10]) >= ex_input1[11:0];
assign jud_12_9 = ((def_12_8<<1'd1) | ex_input0[9]) >= ex_input1[11:0];
assign jud_12_10 = ((def_12_9<<1'd1) | ex_input0[8]) >= ex_input1[11:0];
assign jud_12_11 = ((def_12_10<<1'd1) | ex_input0[7]) >= ex_input1[11:0];
assign jud_12_12 = ((def_12_11<<1'd1) | ex_input0[6]) >= ex_input1[11:0];
assign jud_12_13 = ((def_12_12<<1'd1) | ex_input0[5]) >= ex_input1[11:0];
assign jud_12_14 = ((def_12_13<<1'd1) | ex_input0[4]) >= ex_input1[11:0];
assign jud_12_15 = ((def_12_14<<1'd1) | ex_input0[3]) >= ex_input1[11:0];
assign jud_12_16 = ((def_12_15<<1'd1) | ex_input0[2]) >= ex_input1[11:0];
assign jud_12_17 = ((def_12_16<<1'd1) | ex_input0[1]) >= ex_input1[11:0];
assign jud_12_18 = ((def_12_17<<1'd1) | ex_input0[0]) >= ex_input1[11:0];

assign def_12_0 = ex_input0[29:18] - (ex_input1[11:0] & {5'd12{jud_12_0}});
assign def_12_1 = ((def_12_0<<1'd1) | ex_input0[17]) - (ex_input1[11:0] & {5'd12{jud_12_1}});
assign def_12_2 = ((def_12_1<<1'd1) | ex_input0[16]) - (ex_input1[11:0] & {5'd12{jud_12_2}});
assign def_12_3 = ((def_12_2<<1'd1) | ex_input0[15]) - (ex_input1[11:0] & {5'd12{jud_12_3}});
assign def_12_4 = ((def_12_3<<1'd1) | ex_input0[14]) - (ex_input1[11:0] & {5'd12{jud_12_4}});
assign def_12_5 = ((def_12_4<<1'd1) | ex_input0[13]) - (ex_input1[11:0] & {5'd12{jud_12_5}});
assign def_12_6 = ((def_12_5<<1'd1) | ex_input0[12]) - (ex_input1[11:0] & {5'd12{jud_12_6}});
assign def_12_7 = ((def_12_6<<1'd1) | ex_input0[11]) - (ex_input1[11:0] & {5'd12{jud_12_7}});
assign def_12_8 = ((def_12_7<<1'd1) | ex_input0[10]) - (ex_input1[11:0] & {5'd12{jud_12_8}});
assign def_12_9 = ((def_12_8<<1'd1) | ex_input0[9]) - (ex_input1[11:0] & {5'd12{jud_12_9}});
assign def_12_10 = ((def_12_9<<1'd1) | ex_input0[8]) - (ex_input1[11:0] & {5'd12{jud_12_10}});
assign def_12_11 = ((def_12_10<<1'd1) | ex_input0[7]) - (ex_input1[11:0] & {5'd12{jud_12_11}});
assign def_12_12 = ((def_12_11<<1'd1) | ex_input0[6]) - (ex_input1[11:0] & {5'd12{jud_12_12}});
assign def_12_13 = ((def_12_12<<1'd1) | ex_input0[5]) - (ex_input1[11:0] & {5'd12{jud_12_13}});
assign def_12_14 = ((def_12_13<<1'd1) | ex_input0[4]) - (ex_input1[11:0] & {5'd12{jud_12_14}});
assign def_12_15 = ((def_12_14<<1'd1) | ex_input0[3]) - (ex_input1[11:0] & {5'd12{jud_12_15}});
assign def_12_16 = ((def_12_15<<1'd1) | ex_input0[2]) - (ex_input1[11:0] & {5'd12{jud_12_16}});
assign def_12_17 = ((def_12_16<<1'd1) | ex_input0[1]) - (ex_input1[11:0] & {5'd12{jud_12_17}});
assign def_12_18 = ((def_12_17<<1'd1) | ex_input0[0]) - (ex_input1[11:0] & {5'd12{jud_12_18}});

assign ans_12[29] = 1'd0;
assign ans_12[28] = 1'd0;
assign ans_12[27] = 1'd0;
assign ans_12[26] = 1'd0;
assign ans_12[25] = 1'd0;
assign ans_12[24] = 1'd0;
assign ans_12[23] = 1'd0;
assign ans_12[22] = 1'd0;
assign ans_12[21] = 1'd0;
assign ans_12[20] = 1'd0;
assign ans_12[19] = 1'd0;
assign ans_12[18] = jud_12_0;
assign ans_12[17] = jud_12_1;
assign ans_12[16] = jud_12_2;
assign ans_12[15] = jud_12_3;
assign ans_12[14] = jud_12_4;
assign ans_12[13] = jud_12_5;
assign ans_12[12] = jud_12_6;
assign ans_12[11] = jud_12_7;
assign ans_12[10] = jud_12_8;
assign ans_12[9] = jud_12_9;
assign ans_12[8] = jud_12_10;
assign ans_12[7] = jud_12_11;
assign ans_12[6] = jud_12_12;
assign ans_12[5] = jud_12_13;
assign ans_12[4] = jud_12_14;
assign ans_12[3] = jud_12_15;
assign ans_12[2] = jud_12_16;
assign ans_12[1] = jud_12_17;
assign ans_12[0] = jud_12_18;

// 11bit /////////////////////////////////////////////////////////////////////////////
assign jud_11_0 = ex_input0[29:19] >= ex_input1[10:0];
assign jud_11_1 = ((def_11_0<<1'd1) | ex_input0[18]) >= ex_input1[10:0];
assign jud_11_2 = ((def_11_1<<1'd1) | ex_input0[17]) >= ex_input1[10:0];
assign jud_11_3 = ((def_11_2<<1'd1) | ex_input0[16]) >= ex_input1[10:0];
assign jud_11_4 = ((def_11_3<<1'd1) | ex_input0[15]) >= ex_input1[10:0];
assign jud_11_5 = ((def_11_4<<1'd1) | ex_input0[14]) >= ex_input1[10:0];
assign jud_11_6 = ((def_11_5<<1'd1) | ex_input0[13]) >= ex_input1[10:0];
assign jud_11_7 = ((def_11_6<<1'd1) | ex_input0[12]) >= ex_input1[10:0];
assign jud_11_8 = ((def_11_7<<1'd1) | ex_input0[11]) >= ex_input1[10:0];
assign jud_11_9 = ((def_11_8<<1'd1) | ex_input0[10]) >= ex_input1[10:0];
assign jud_11_10 = ((def_11_9<<1'd1) | ex_input0[9]) >= ex_input1[10:0];
assign jud_11_11 = ((def_11_10<<1'd1) | ex_input0[8]) >= ex_input1[10:0];
assign jud_11_12 = ((def_11_11<<1'd1) | ex_input0[7]) >= ex_input1[10:0];
assign jud_11_13 = ((def_11_12<<1'd1) | ex_input0[6]) >= ex_input1[10:0];
assign jud_11_14 = ((def_11_13<<1'd1) | ex_input0[5]) >= ex_input1[10:0];
assign jud_11_15 = ((def_11_14<<1'd1) | ex_input0[4]) >= ex_input1[10:0];
assign jud_11_16 = ((def_11_15<<1'd1) | ex_input0[3]) >= ex_input1[10:0];
assign jud_11_17 = ((def_11_16<<1'd1) | ex_input0[2]) >= ex_input1[10:0];
assign jud_11_18 = ((def_11_17<<1'd1) | ex_input0[1]) >= ex_input1[10:0];
assign jud_11_19 = ((def_11_18<<1'd1) | ex_input0[0]) >= ex_input1[10:0];

assign def_11_0 = ex_input0[29:19] - (ex_input1[10:0] & {5'd11{jud_11_0}});
assign def_11_1 = ((def_11_0<<1'd1) | ex_input0[18]) - (ex_input1[10:0] & {5'd11{jud_11_1}});
assign def_11_2 = ((def_11_1<<1'd1) | ex_input0[17]) - (ex_input1[10:0] & {5'd11{jud_11_2}});
assign def_11_3 = ((def_11_2<<1'd1) | ex_input0[16]) - (ex_input1[10:0] & {5'd11{jud_11_3}});
assign def_11_4 = ((def_11_3<<1'd1) | ex_input0[15]) - (ex_input1[10:0] & {5'd11{jud_11_4}});
assign def_11_5 = ((def_11_4<<1'd1) | ex_input0[14]) - (ex_input1[10:0] & {5'd11{jud_11_5}});
assign def_11_6 = ((def_11_5<<1'd1) | ex_input0[13]) - (ex_input1[10:0] & {5'd11{jud_11_6}});
assign def_11_7 = ((def_11_6<<1'd1) | ex_input0[12]) - (ex_input1[10:0] & {5'd11{jud_11_7}});
assign def_11_8 = ((def_11_7<<1'd1) | ex_input0[11]) - (ex_input1[10:0] & {5'd11{jud_11_8}});
assign def_11_9 = ((def_11_8<<1'd1) | ex_input0[10]) - (ex_input1[10:0] & {5'd11{jud_11_9}});
assign def_11_10 = ((def_11_9<<1'd1) | ex_input0[9]) - (ex_input1[10:0] & {5'd11{jud_11_10}});
assign def_11_11 = ((def_11_10<<1'd1) | ex_input0[8]) - (ex_input1[10:0] & {5'd11{jud_11_11}});
assign def_11_12 = ((def_11_11<<1'd1) | ex_input0[7]) - (ex_input1[10:0] & {5'd11{jud_11_12}});
assign def_11_13 = ((def_11_12<<1'd1) | ex_input0[6]) - (ex_input1[10:0] & {5'd11{jud_11_13}});
assign def_11_14 = ((def_11_13<<1'd1) | ex_input0[5]) - (ex_input1[10:0] & {5'd11{jud_11_14}});
assign def_11_15 = ((def_11_14<<1'd1) | ex_input0[4]) - (ex_input1[10:0] & {5'd11{jud_11_15}});
assign def_11_16 = ((def_11_15<<1'd1) | ex_input0[3]) - (ex_input1[10:0] & {5'd11{jud_11_16}});
assign def_11_17 = ((def_11_16<<1'd1) | ex_input0[2]) - (ex_input1[10:0] & {5'd11{jud_11_17}});
assign def_11_18 = ((def_11_17<<1'd1) | ex_input0[1]) - (ex_input1[10:0] & {5'd11{jud_11_18}});
assign def_11_19 = ((def_11_18<<1'd1) | ex_input0[0]) - (ex_input1[10:0] & {5'd11{jud_11_19}});

assign ans_11[29] = 1'd0;
assign ans_11[28] = 1'd0;
assign ans_11[27] = 1'd0;
assign ans_11[26] = 1'd0;
assign ans_11[25] = 1'd0;
assign ans_11[24] = 1'd0;
assign ans_11[23] = 1'd0;
assign ans_11[22] = 1'd0;
assign ans_11[21] = 1'd0;
assign ans_11[20] = 1'd0;
assign ans_11[19] = jud_11_0;
assign ans_11[18] = jud_11_1;
assign ans_11[17] = jud_11_2;
assign ans_11[16] = jud_11_3;
assign ans_11[15] = jud_11_4;
assign ans_11[14] = jud_11_5;
assign ans_11[13] = jud_11_6;
assign ans_11[12] = jud_11_7;
assign ans_11[11] = jud_11_8;
assign ans_11[10] = jud_11_9;
assign ans_11[9] = jud_11_10;
assign ans_11[8] = jud_11_11;
assign ans_11[7] = jud_11_12;
assign ans_11[6] = jud_11_13;
assign ans_11[5] = jud_11_14;
assign ans_11[4] = jud_11_15;
assign ans_11[3] = jud_11_16;
assign ans_11[2] = jud_11_17;
assign ans_11[1] = jud_11_18;
assign ans_11[0] = jud_11_19;

// 10bit /////////////////////////////////////////////////////////////////////////////
assign jud_10_0 = ex_input0[29:20] >= ex_input1[9:0];
assign jud_10_1 = ((def_10_0<<1'd1) | ex_input0[19]) >= ex_input1[9:0];
assign jud_10_2 = ((def_10_1<<1'd1) | ex_input0[18]) >= ex_input1[9:0];
assign jud_10_3 = ((def_10_2<<1'd1) | ex_input0[17]) >= ex_input1[9:0];
assign jud_10_4 = ((def_10_3<<1'd1) | ex_input0[16]) >= ex_input1[9:0];
assign jud_10_5 = ((def_10_4<<1'd1) | ex_input0[15]) >= ex_input1[9:0];
assign jud_10_6 = ((def_10_5<<1'd1) | ex_input0[14]) >= ex_input1[9:0];
assign jud_10_7 = ((def_10_6<<1'd1) | ex_input0[13]) >= ex_input1[9:0];
assign jud_10_8 = ((def_10_7<<1'd1) | ex_input0[12]) >= ex_input1[9:0];
assign jud_10_9 = ((def_10_8<<1'd1) | ex_input0[11]) >= ex_input1[9:0];
assign jud_10_10 = ((def_10_9<<1'd1) | ex_input0[10]) >= ex_input1[9:0];
assign jud_10_11 = ((def_10_10<<1'd1) | ex_input0[9]) >= ex_input1[9:0];
assign jud_10_12 = ((def_10_11<<1'd1) | ex_input0[8]) >= ex_input1[9:0];
assign jud_10_13 = ((def_10_12<<1'd1) | ex_input0[7]) >= ex_input1[9:0];
assign jud_10_14 = ((def_10_13<<1'd1) | ex_input0[6]) >= ex_input1[9:0];
assign jud_10_15 = ((def_10_14<<1'd1) | ex_input0[5]) >= ex_input1[9:0];
assign jud_10_16 = ((def_10_15<<1'd1) | ex_input0[4]) >= ex_input1[9:0];
assign jud_10_17 = ((def_10_16<<1'd1) | ex_input0[3]) >= ex_input1[9:0];
assign jud_10_18 = ((def_10_17<<1'd1) | ex_input0[2]) >= ex_input1[9:0];
assign jud_10_19 = ((def_10_18<<1'd1) | ex_input0[1]) >= ex_input1[9:0];
assign jud_10_20 = ((def_10_19<<1'd1) | ex_input0[0]) >= ex_input1[9:0];

assign def_10_0 = ex_input0[29:20] - (ex_input1[9:0] & {5'd10{jud_10_0}});
assign def_10_1 = ((def_10_0<<1'd1) | ex_input0[19]) - (ex_input1[9:0] & {5'd10{jud_10_1}});
assign def_10_2 = ((def_10_1<<1'd1) | ex_input0[18]) - (ex_input1[9:0] & {5'd10{jud_10_2}});
assign def_10_3 = ((def_10_2<<1'd1) | ex_input0[17]) - (ex_input1[9:0] & {5'd10{jud_10_3}});
assign def_10_4 = ((def_10_3<<1'd1) | ex_input0[16]) - (ex_input1[9:0] & {5'd10{jud_10_4}});
assign def_10_5 = ((def_10_4<<1'd1) | ex_input0[15]) - (ex_input1[9:0] & {5'd10{jud_10_5}});
assign def_10_6 = ((def_10_5<<1'd1) | ex_input0[14]) - (ex_input1[9:0] & {5'd10{jud_10_6}});
assign def_10_7 = ((def_10_6<<1'd1) | ex_input0[13]) - (ex_input1[9:0] & {5'd10{jud_10_7}});
assign def_10_8 = ((def_10_7<<1'd1) | ex_input0[12]) - (ex_input1[9:0] & {5'd10{jud_10_8}});
assign def_10_9 = ((def_10_8<<1'd1) | ex_input0[11]) - (ex_input1[9:0] & {5'd10{jud_10_9}});
assign def_10_10 = ((def_10_9<<1'd1) | ex_input0[10]) - (ex_input1[9:0] & {5'd10{jud_10_10}});
assign def_10_11 = ((def_10_10<<1'd1) | ex_input0[9]) - (ex_input1[9:0] & {5'd10{jud_10_11}});
assign def_10_12 = ((def_10_11<<1'd1) | ex_input0[8]) - (ex_input1[9:0] & {5'd10{jud_10_12}});
assign def_10_13 = ((def_10_12<<1'd1) | ex_input0[7]) - (ex_input1[9:0] & {5'd10{jud_10_13}});
assign def_10_14 = ((def_10_13<<1'd1) | ex_input0[6]) - (ex_input1[9:0] & {5'd10{jud_10_14}});
assign def_10_15 = ((def_10_14<<1'd1) | ex_input0[5]) - (ex_input1[9:0] & {5'd10{jud_10_15}});
assign def_10_16 = ((def_10_15<<1'd1) | ex_input0[4]) - (ex_input1[9:0] & {5'd10{jud_10_16}});
assign def_10_17 = ((def_10_16<<1'd1) | ex_input0[3]) - (ex_input1[9:0] & {5'd10{jud_10_17}});
assign def_10_18 = ((def_10_17<<1'd1) | ex_input0[2]) - (ex_input1[9:0] & {5'd10{jud_10_18}});
assign def_10_19 = ((def_10_18<<1'd1) | ex_input0[1]) - (ex_input1[9:0] & {5'd10{jud_10_19}});
assign def_10_20 = ((def_10_19<<1'd1) | ex_input0[0]) - (ex_input1[9:0] & {5'd10{jud_10_20}});

assign ans_10[29] = 1'd0;
assign ans_10[28] = 1'd0;
assign ans_10[27] = 1'd0;
assign ans_10[26] = 1'd0;
assign ans_10[25] = 1'd0;
assign ans_10[24] = 1'd0;
assign ans_10[23] = 1'd0;
assign ans_10[22] = 1'd0;
assign ans_10[21] = 1'd0;
assign ans_10[20] = jud_10_0;
assign ans_10[19] = jud_10_1;
assign ans_10[18] = jud_10_2;
assign ans_10[17] = jud_10_3;
assign ans_10[16] = jud_10_4;
assign ans_10[15] = jud_10_5;
assign ans_10[14] = jud_10_6;
assign ans_10[13] = jud_10_7;
assign ans_10[12] = jud_10_8;
assign ans_10[11] = jud_10_9;
assign ans_10[10] = jud_10_10;
assign ans_10[9] = jud_10_11;
assign ans_10[8] = jud_10_12;
assign ans_10[7] = jud_10_13;
assign ans_10[6] = jud_10_14;
assign ans_10[5] = jud_10_15;
assign ans_10[4] = jud_10_16;
assign ans_10[3] = jud_10_17;
assign ans_10[2] = jud_10_18;
assign ans_10[1] = jud_10_19;
assign ans_10[0] = jud_10_20;

//  9bit /////////////////////////////////////////////////////////////////////////////
assign jud_9_0 = ex_input0[29:21] >= ex_input1[8:0];
assign jud_9_1 = ((def_9_0<<1'd1) | ex_input0[20]) >= ex_input1[8:0];
assign jud_9_2 = ((def_9_1<<1'd1) | ex_input0[19]) >= ex_input1[8:0];
assign jud_9_3 = ((def_9_2<<1'd1) | ex_input0[18]) >= ex_input1[8:0];
assign jud_9_4 = ((def_9_3<<1'd1) | ex_input0[17]) >= ex_input1[8:0];
assign jud_9_5 = ((def_9_4<<1'd1) | ex_input0[16]) >= ex_input1[8:0];
assign jud_9_6 = ((def_9_5<<1'd1) | ex_input0[15]) >= ex_input1[8:0];
assign jud_9_7 = ((def_9_6<<1'd1) | ex_input0[14]) >= ex_input1[8:0];
assign jud_9_8 = ((def_9_7<<1'd1) | ex_input0[13]) >= ex_input1[8:0];
assign jud_9_9 = ((def_9_8<<1'd1) | ex_input0[12]) >= ex_input1[8:0];
assign jud_9_10 = ((def_9_9<<1'd1) | ex_input0[11]) >= ex_input1[8:0];
assign jud_9_11 = ((def_9_10<<1'd1) | ex_input0[10]) >= ex_input1[8:0];
assign jud_9_12 = ((def_9_11<<1'd1) | ex_input0[9]) >= ex_input1[8:0];
assign jud_9_13 = ((def_9_12<<1'd1) | ex_input0[8]) >= ex_input1[8:0];
assign jud_9_14 = ((def_9_13<<1'd1) | ex_input0[7]) >= ex_input1[8:0];
assign jud_9_15 = ((def_9_14<<1'd1) | ex_input0[6]) >= ex_input1[8:0];
assign jud_9_16 = ((def_9_15<<1'd1) | ex_input0[5]) >= ex_input1[8:0];
assign jud_9_17 = ((def_9_16<<1'd1) | ex_input0[4]) >= ex_input1[8:0];
assign jud_9_18 = ((def_9_17<<1'd1) | ex_input0[3]) >= ex_input1[8:0];
assign jud_9_19 = ((def_9_18<<1'd1) | ex_input0[2]) >= ex_input1[8:0];
assign jud_9_20 = ((def_9_19<<1'd1) | ex_input0[1]) >= ex_input1[8:0];
assign jud_9_21 = ((def_9_20<<1'd1) | ex_input0[0]) >= ex_input1[8:0];

assign def_9_0 = ex_input0[29:21] - (ex_input1[8:0] & {5'd9{jud_9_0}});
assign def_9_1 = ((def_9_0<<1'd1) | ex_input0[20]) - (ex_input1[8:0] & {5'd9{jud_9_1}});
assign def_9_2 = ((def_9_1<<1'd1) | ex_input0[19]) - (ex_input1[8:0] & {5'd9{jud_9_2}});
assign def_9_3 = ((def_9_2<<1'd1) | ex_input0[18]) - (ex_input1[8:0] & {5'd9{jud_9_3}});
assign def_9_4 = ((def_9_3<<1'd1) | ex_input0[17]) - (ex_input1[8:0] & {5'd9{jud_9_4}});
assign def_9_5 = ((def_9_4<<1'd1) | ex_input0[16]) - (ex_input1[8:0] & {5'd9{jud_9_5}});
assign def_9_6 = ((def_9_5<<1'd1) | ex_input0[15]) - (ex_input1[8:0] & {5'd9{jud_9_6}});
assign def_9_7 = ((def_9_6<<1'd1) | ex_input0[14]) - (ex_input1[8:0] & {5'd9{jud_9_7}});
assign def_9_8 = ((def_9_7<<1'd1) | ex_input0[13]) - (ex_input1[8:0] & {5'd9{jud_9_8}});
assign def_9_9 = ((def_9_8<<1'd1) | ex_input0[12]) - (ex_input1[8:0] & {5'd9{jud_9_9}});
assign def_9_10 = ((def_9_9<<1'd1) | ex_input0[11]) - (ex_input1[8:0] & {5'd9{jud_9_10}});
assign def_9_11 = ((def_9_10<<1'd1) | ex_input0[10]) - (ex_input1[8:0] & {5'd9{jud_9_11}});
assign def_9_12 = ((def_9_11<<1'd1) | ex_input0[9]) - (ex_input1[8:0] & {5'd9{jud_9_12}});
assign def_9_13 = ((def_9_12<<1'd1) | ex_input0[8]) - (ex_input1[8:0] & {5'd9{jud_9_13}});
assign def_9_14 = ((def_9_13<<1'd1) | ex_input0[7]) - (ex_input1[8:0] & {5'd9{jud_9_14}});
assign def_9_15 = ((def_9_14<<1'd1) | ex_input0[6]) - (ex_input1[8:0] & {5'd9{jud_9_15}});
assign def_9_16 = ((def_9_15<<1'd1) | ex_input0[5]) - (ex_input1[8:0] & {5'd9{jud_9_16}});
assign def_9_17 = ((def_9_16<<1'd1) | ex_input0[4]) - (ex_input1[8:0] & {5'd9{jud_9_17}});
assign def_9_18 = ((def_9_17<<1'd1) | ex_input0[3]) - (ex_input1[8:0] & {5'd9{jud_9_18}});
assign def_9_19 = ((def_9_18<<1'd1) | ex_input0[2]) - (ex_input1[8:0] & {5'd9{jud_9_19}});
assign def_9_20 = ((def_9_19<<1'd1) | ex_input0[1]) - (ex_input1[8:0] & {5'd9{jud_9_20}});
assign def_9_21 = ((def_9_20<<1'd1) | ex_input0[0]) - (ex_input1[8:0] & {5'd9{jud_9_21}});

assign ans_9[29] = 1'd0;
assign ans_9[28] = 1'd0;
assign ans_9[27] = 1'd0;
assign ans_9[26] = 1'd0;
assign ans_9[25] = 1'd0;
assign ans_9[24] = 1'd0;
assign ans_9[23] = 1'd0;
assign ans_9[22] = 1'd0;
assign ans_9[21] = jud_9_0;
assign ans_9[20] = jud_9_1;
assign ans_9[19] = jud_9_2;
assign ans_9[18] = jud_9_3;
assign ans_9[17] = jud_9_4;
assign ans_9[16] = jud_9_5;
assign ans_9[15] = jud_9_6;
assign ans_9[14] = jud_9_7;
assign ans_9[13] = jud_9_8;
assign ans_9[12] = jud_9_9;
assign ans_9[11] = jud_9_10;
assign ans_9[10] = jud_9_11;
assign ans_9[9] = jud_9_12;
assign ans_9[8] = jud_9_13;
assign ans_9[7] = jud_9_14;
assign ans_9[6] = jud_9_15;
assign ans_9[5] = jud_9_16;
assign ans_9[4] = jud_9_17;
assign ans_9[3] = jud_9_18;
assign ans_9[2] = jud_9_19;
assign ans_9[1] = jud_9_20;
assign ans_9[0] = jud_9_21;

//  8bit /////////////////////////////////////////////////////////////////////////////
assign jud_8_0 = ex_input0[29:22] >= ex_input1[7:0];
assign jud_8_1 = ((def_8_0<<1'd1) | ex_input0[21]) >= ex_input1[7:0];
assign jud_8_2 = ((def_8_1<<1'd1) | ex_input0[20]) >= ex_input1[7:0];
assign jud_8_3 = ((def_8_2<<1'd1) | ex_input0[19]) >= ex_input1[7:0];
assign jud_8_4 = ((def_8_3<<1'd1) | ex_input0[18]) >= ex_input1[7:0];
assign jud_8_5 = ((def_8_4<<1'd1) | ex_input0[17]) >= ex_input1[7:0];
assign jud_8_6 = ((def_8_5<<1'd1) | ex_input0[16]) >= ex_input1[7:0];
assign jud_8_7 = ((def_8_6<<1'd1) | ex_input0[15]) >= ex_input1[7:0];
assign jud_8_8 = ((def_8_7<<1'd1) | ex_input0[14]) >= ex_input1[7:0];
assign jud_8_9 = ((def_8_8<<1'd1) | ex_input0[13]) >= ex_input1[7:0];
assign jud_8_10 = ((def_8_9<<1'd1) | ex_input0[12]) >= ex_input1[7:0];
assign jud_8_11 = ((def_8_10<<1'd1) | ex_input0[11]) >= ex_input1[7:0];
assign jud_8_12 = ((def_8_11<<1'd1) | ex_input0[10]) >= ex_input1[7:0];
assign jud_8_13 = ((def_8_12<<1'd1) | ex_input0[9]) >= ex_input1[7:0];
assign jud_8_14 = ((def_8_13<<1'd1) | ex_input0[8]) >= ex_input1[7:0];
assign jud_8_15 = ((def_8_14<<1'd1) | ex_input0[7]) >= ex_input1[7:0];
assign jud_8_16 = ((def_8_15<<1'd1) | ex_input0[6]) >= ex_input1[7:0];
assign jud_8_17 = ((def_8_16<<1'd1) | ex_input0[5]) >= ex_input1[7:0];
assign jud_8_18 = ((def_8_17<<1'd1) | ex_input0[4]) >= ex_input1[7:0];
assign jud_8_19 = ((def_8_18<<1'd1) | ex_input0[3]) >= ex_input1[7:0];
assign jud_8_20 = ((def_8_19<<1'd1) | ex_input0[2]) >= ex_input1[7:0];
assign jud_8_21 = ((def_8_20<<1'd1) | ex_input0[1]) >= ex_input1[7:0];
assign jud_8_22 = ((def_8_21<<1'd1) | ex_input0[0]) >= ex_input1[7:0];

assign def_8_0 = ex_input0[29:22] - (ex_input1[7:0] & {5'd8{jud_8_0}});
assign def_8_1 = ((def_8_0<<1'd1) | ex_input0[21]) - (ex_input1[7:0] & {5'd8{jud_8_1}});
assign def_8_2 = ((def_8_1<<1'd1) | ex_input0[20]) - (ex_input1[7:0] & {5'd8{jud_8_2}});
assign def_8_3 = ((def_8_2<<1'd1) | ex_input0[19]) - (ex_input1[7:0] & {5'd8{jud_8_3}});
assign def_8_4 = ((def_8_3<<1'd1) | ex_input0[18]) - (ex_input1[7:0] & {5'd8{jud_8_4}});
assign def_8_5 = ((def_8_4<<1'd1) | ex_input0[17]) - (ex_input1[7:0] & {5'd8{jud_8_5}});
assign def_8_6 = ((def_8_5<<1'd1) | ex_input0[16]) - (ex_input1[7:0] & {5'd8{jud_8_6}});
assign def_8_7 = ((def_8_6<<1'd1) | ex_input0[15]) - (ex_input1[7:0] & {5'd8{jud_8_7}});
assign def_8_8 = ((def_8_7<<1'd1) | ex_input0[14]) - (ex_input1[7:0] & {5'd8{jud_8_8}});
assign def_8_9 = ((def_8_8<<1'd1) | ex_input0[13]) - (ex_input1[7:0] & {5'd8{jud_8_9}});
assign def_8_10 = ((def_8_9<<1'd1) | ex_input0[12]) - (ex_input1[7:0] & {5'd8{jud_8_10}});
assign def_8_11 = ((def_8_10<<1'd1) | ex_input0[11]) - (ex_input1[7:0] & {5'd8{jud_8_11}});
assign def_8_12 = ((def_8_11<<1'd1) | ex_input0[10]) - (ex_input1[7:0] & {5'd8{jud_8_12}});
assign def_8_13 = ((def_8_12<<1'd1) | ex_input0[9]) - (ex_input1[7:0] & {5'd8{jud_8_13}});
assign def_8_14 = ((def_8_13<<1'd1) | ex_input0[8]) - (ex_input1[7:0] & {5'd8{jud_8_14}});
assign def_8_15 = ((def_8_14<<1'd1) | ex_input0[7]) - (ex_input1[7:0] & {5'd8{jud_8_15}});
assign def_8_16 = ((def_8_15<<1'd1) | ex_input0[6]) - (ex_input1[7:0] & {5'd8{jud_8_16}});
assign def_8_17 = ((def_8_16<<1'd1) | ex_input0[5]) - (ex_input1[7:0] & {5'd8{jud_8_17}});
assign def_8_18 = ((def_8_17<<1'd1) | ex_input0[4]) - (ex_input1[7:0] & {5'd8{jud_8_18}});
assign def_8_19 = ((def_8_18<<1'd1) | ex_input0[3]) - (ex_input1[7:0] & {5'd8{jud_8_19}});
assign def_8_20 = ((def_8_19<<1'd1) | ex_input0[2]) - (ex_input1[7:0] & {5'd8{jud_8_20}});
assign def_8_21 = ((def_8_20<<1'd1) | ex_input0[1]) - (ex_input1[7:0] & {5'd8{jud_8_21}});
assign def_8_22 = ((def_8_21<<1'd1) | ex_input0[0]) - (ex_input1[7:0] & {5'd8{jud_8_22}});

assign ans_8[29] = 1'd0;
assign ans_8[28] = 1'd0;
assign ans_8[27] = 1'd0;
assign ans_8[26] = 1'd0;
assign ans_8[25] = 1'd0;
assign ans_8[24] = 1'd0;
assign ans_8[23] = 1'd0;
assign ans_8[22] = jud_8_0;
assign ans_8[21] = jud_8_1;
assign ans_8[20] = jud_8_2;
assign ans_8[19] = jud_8_3;
assign ans_8[18] = jud_8_4;
assign ans_8[17] = jud_8_5;
assign ans_8[16] = jud_8_6;
assign ans_8[15] = jud_8_7;
assign ans_8[14] = jud_8_8;
assign ans_8[13] = jud_8_9;
assign ans_8[12] = jud_8_10;
assign ans_8[11] = jud_8_11;
assign ans_8[10] = jud_8_12;
assign ans_8[9] = jud_8_13;
assign ans_8[8] = jud_8_14;
assign ans_8[7] = jud_8_15;
assign ans_8[6] = jud_8_16;
assign ans_8[5] = jud_8_17;
assign ans_8[4] = jud_8_18;
assign ans_8[3] = jud_8_19;
assign ans_8[2] = jud_8_20;
assign ans_8[1] = jud_8_21;
assign ans_8[0] = jud_8_22;

//  7bit /////////////////////////////////////////////////////////////////////////////
assign jud_7_0 = ex_input0[29:23] >= ex_input1[6:0];
assign jud_7_1 = ((def_7_0<<1'd1) | ex_input0[22]) >= ex_input1[6:0];
assign jud_7_2 = ((def_7_1<<1'd1) | ex_input0[21]) >= ex_input1[6:0];
assign jud_7_3 = ((def_7_2<<1'd1) | ex_input0[20]) >= ex_input1[6:0];
assign jud_7_4 = ((def_7_3<<1'd1) | ex_input0[19]) >= ex_input1[6:0];
assign jud_7_5 = ((def_7_4<<1'd1) | ex_input0[18]) >= ex_input1[6:0];
assign jud_7_6 = ((def_7_5<<1'd1) | ex_input0[17]) >= ex_input1[6:0];
assign jud_7_7 = ((def_7_6<<1'd1) | ex_input0[16]) >= ex_input1[6:0];
assign jud_7_8 = ((def_7_7<<1'd1) | ex_input0[15]) >= ex_input1[6:0];
assign jud_7_9 = ((def_7_8<<1'd1) | ex_input0[14]) >= ex_input1[6:0];
assign jud_7_10 = ((def_7_9<<1'd1) | ex_input0[13]) >= ex_input1[6:0];
assign jud_7_11 = ((def_7_10<<1'd1) | ex_input0[12]) >= ex_input1[6:0];
assign jud_7_12 = ((def_7_11<<1'd1) | ex_input0[11]) >= ex_input1[6:0];
assign jud_7_13 = ((def_7_12<<1'd1) | ex_input0[10]) >= ex_input1[6:0];
assign jud_7_14 = ((def_7_13<<1'd1) | ex_input0[9]) >= ex_input1[6:0];
assign jud_7_15 = ((def_7_14<<1'd1) | ex_input0[8]) >= ex_input1[6:0];
assign jud_7_16 = ((def_7_15<<1'd1) | ex_input0[7]) >= ex_input1[6:0];
assign jud_7_17 = ((def_7_16<<1'd1) | ex_input0[6]) >= ex_input1[6:0];
assign jud_7_18 = ((def_7_17<<1'd1) | ex_input0[5]) >= ex_input1[6:0];
assign jud_7_19 = ((def_7_18<<1'd1) | ex_input0[4]) >= ex_input1[6:0];
assign jud_7_20 = ((def_7_19<<1'd1) | ex_input0[3]) >= ex_input1[6:0];
assign jud_7_21 = ((def_7_20<<1'd1) | ex_input0[2]) >= ex_input1[6:0];
assign jud_7_22 = ((def_7_21<<1'd1) | ex_input0[1]) >= ex_input1[6:0];
assign jud_7_23 = ((def_7_22<<1'd1) | ex_input0[0]) >= ex_input1[6:0];

assign def_7_0 = ex_input0[29:23] - (ex_input1[6:0] & {5'd7{jud_7_0}});
assign def_7_1 = ((def_7_0<<1'd1) | ex_input0[22]) - (ex_input1[6:0] & {5'd7{jud_7_1}});
assign def_7_2 = ((def_7_1<<1'd1) | ex_input0[21]) - (ex_input1[6:0] & {5'd7{jud_7_2}});
assign def_7_3 = ((def_7_2<<1'd1) | ex_input0[20]) - (ex_input1[6:0] & {5'd7{jud_7_3}});
assign def_7_4 = ((def_7_3<<1'd1) | ex_input0[19]) - (ex_input1[6:0] & {5'd7{jud_7_4}});
assign def_7_5 = ((def_7_4<<1'd1) | ex_input0[18]) - (ex_input1[6:0] & {5'd7{jud_7_5}});
assign def_7_6 = ((def_7_5<<1'd1) | ex_input0[17]) - (ex_input1[6:0] & {5'd7{jud_7_6}});
assign def_7_7 = ((def_7_6<<1'd1) | ex_input0[16]) - (ex_input1[6:0] & {5'd7{jud_7_7}});
assign def_7_8 = ((def_7_7<<1'd1) | ex_input0[15]) - (ex_input1[6:0] & {5'd7{jud_7_8}});
assign def_7_9 = ((def_7_8<<1'd1) | ex_input0[14]) - (ex_input1[6:0] & {5'd7{jud_7_9}});
assign def_7_10 = ((def_7_9<<1'd1) | ex_input0[13]) - (ex_input1[6:0] & {5'd7{jud_7_10}});
assign def_7_11 = ((def_7_10<<1'd1) | ex_input0[12]) - (ex_input1[6:0] & {5'd7{jud_7_11}});
assign def_7_12 = ((def_7_11<<1'd1) | ex_input0[11]) - (ex_input1[6:0] & {5'd7{jud_7_12}});
assign def_7_13 = ((def_7_12<<1'd1) | ex_input0[10]) - (ex_input1[6:0] & {5'd7{jud_7_13}});
assign def_7_14 = ((def_7_13<<1'd1) | ex_input0[9]) - (ex_input1[6:0] & {5'd7{jud_7_14}});
assign def_7_15 = ((def_7_14<<1'd1) | ex_input0[8]) - (ex_input1[6:0] & {5'd7{jud_7_15}});
assign def_7_16 = ((def_7_15<<1'd1) | ex_input0[7]) - (ex_input1[6:0] & {5'd7{jud_7_16}});
assign def_7_17 = ((def_7_16<<1'd1) | ex_input0[6]) - (ex_input1[6:0] & {5'd7{jud_7_17}});
assign def_7_18 = ((def_7_17<<1'd1) | ex_input0[5]) - (ex_input1[6:0] & {5'd7{jud_7_18}});
assign def_7_19 = ((def_7_18<<1'd1) | ex_input0[4]) - (ex_input1[6:0] & {5'd7{jud_7_19}});
assign def_7_20 = ((def_7_19<<1'd1) | ex_input0[3]) - (ex_input1[6:0] & {5'd7{jud_7_20}});
assign def_7_21 = ((def_7_20<<1'd1) | ex_input0[2]) - (ex_input1[6:0] & {5'd7{jud_7_21}});
assign def_7_22 = ((def_7_21<<1'd1) | ex_input0[1]) - (ex_input1[6:0] & {5'd7{jud_7_22}});
assign def_7_23 = ((def_7_22<<1'd1) | ex_input0[0]) - (ex_input1[6:0] & {5'd7{jud_7_23}});

assign ans_7[29] = 1'd0;
assign ans_7[28] = 1'd0;
assign ans_7[27] = 1'd0;
assign ans_7[26] = 1'd0;
assign ans_7[25] = 1'd0;
assign ans_7[24] = 1'd0;
assign ans_7[23] = jud_7_0;
assign ans_7[22] = jud_7_1;
assign ans_7[21] = jud_7_2;
assign ans_7[20] = jud_7_3;
assign ans_7[19] = jud_7_4;
assign ans_7[18] = jud_7_5;
assign ans_7[17] = jud_7_6;
assign ans_7[16] = jud_7_7;
assign ans_7[15] = jud_7_8;
assign ans_7[14] = jud_7_9;
assign ans_7[13] = jud_7_10;
assign ans_7[12] = jud_7_11;
assign ans_7[11] = jud_7_12;
assign ans_7[10] = jud_7_13;
assign ans_7[9] = jud_7_14;
assign ans_7[8] = jud_7_15;
assign ans_7[7] = jud_7_16;
assign ans_7[6] = jud_7_17;
assign ans_7[5] = jud_7_18;
assign ans_7[4] = jud_7_19;
assign ans_7[3] = jud_7_20;
assign ans_7[2] = jud_7_21;
assign ans_7[1] = jud_7_22;
assign ans_7[0] = jud_7_23;

//  6bit /////////////////////////////////////////////////////////////////////////////
assign jud_6_0 = ex_input0[29:24] >= ex_input1[5:0];
assign jud_6_1 = ((def_6_0<<1'd1) | ex_input0[23]) >= ex_input1[5:0];
assign jud_6_2 = ((def_6_1<<1'd1) | ex_input0[22]) >= ex_input1[5:0];
assign jud_6_3 = ((def_6_2<<1'd1) | ex_input0[21]) >= ex_input1[5:0];
assign jud_6_4 = ((def_6_3<<1'd1) | ex_input0[20]) >= ex_input1[5:0];
assign jud_6_5 = ((def_6_4<<1'd1) | ex_input0[19]) >= ex_input1[5:0];
assign jud_6_6 = ((def_6_5<<1'd1) | ex_input0[18]) >= ex_input1[5:0];
assign jud_6_7 = ((def_6_6<<1'd1) | ex_input0[17]) >= ex_input1[5:0];
assign jud_6_8 = ((def_6_7<<1'd1) | ex_input0[16]) >= ex_input1[5:0];
assign jud_6_9 = ((def_6_8<<1'd1) | ex_input0[15]) >= ex_input1[5:0];
assign jud_6_10 = ((def_6_9<<1'd1) | ex_input0[14]) >= ex_input1[5:0];
assign jud_6_11 = ((def_6_10<<1'd1) | ex_input0[13]) >= ex_input1[5:0];
assign jud_6_12 = ((def_6_11<<1'd1) | ex_input0[12]) >= ex_input1[5:0];
assign jud_6_13 = ((def_6_12<<1'd1) | ex_input0[11]) >= ex_input1[5:0];
assign jud_6_14 = ((def_6_13<<1'd1) | ex_input0[10]) >= ex_input1[5:0];
assign jud_6_15 = ((def_6_14<<1'd1) | ex_input0[9]) >= ex_input1[5:0];
assign jud_6_16 = ((def_6_15<<1'd1) | ex_input0[8]) >= ex_input1[5:0];
assign jud_6_17 = ((def_6_16<<1'd1) | ex_input0[7]) >= ex_input1[5:0];
assign jud_6_18 = ((def_6_17<<1'd1) | ex_input0[6]) >= ex_input1[5:0];
assign jud_6_19 = ((def_6_18<<1'd1) | ex_input0[5]) >= ex_input1[5:0];
assign jud_6_20 = ((def_6_19<<1'd1) | ex_input0[4]) >= ex_input1[5:0];
assign jud_6_21 = ((def_6_20<<1'd1) | ex_input0[3]) >= ex_input1[5:0];
assign jud_6_22 = ((def_6_21<<1'd1) | ex_input0[2]) >= ex_input1[5:0];
assign jud_6_23 = ((def_6_22<<1'd1) | ex_input0[1]) >= ex_input1[5:0];
assign jud_6_24 = ((def_6_23<<1'd1) | ex_input0[0]) >= ex_input1[5:0];

assign def_6_0 = ex_input0[29:24] - (ex_input1[5:0] & {5'd6{jud_6_0}});
assign def_6_1 = ((def_6_0<<1'd1) | ex_input0[23]) - (ex_input1[5:0] & {5'd6{jud_6_1}});
assign def_6_2 = ((def_6_1<<1'd1) | ex_input0[22]) - (ex_input1[5:0] & {5'd6{jud_6_2}});
assign def_6_3 = ((def_6_2<<1'd1) | ex_input0[21]) - (ex_input1[5:0] & {5'd6{jud_6_3}});
assign def_6_4 = ((def_6_3<<1'd1) | ex_input0[20]) - (ex_input1[5:0] & {5'd6{jud_6_4}});
assign def_6_5 = ((def_6_4<<1'd1) | ex_input0[19]) - (ex_input1[5:0] & {5'd6{jud_6_5}});
assign def_6_6 = ((def_6_5<<1'd1) | ex_input0[18]) - (ex_input1[5:0] & {5'd6{jud_6_6}});
assign def_6_7 = ((def_6_6<<1'd1) | ex_input0[17]) - (ex_input1[5:0] & {5'd6{jud_6_7}});
assign def_6_8 = ((def_6_7<<1'd1) | ex_input0[16]) - (ex_input1[5:0] & {5'd6{jud_6_8}});
assign def_6_9 = ((def_6_8<<1'd1) | ex_input0[15]) - (ex_input1[5:0] & {5'd6{jud_6_9}});
assign def_6_10 = ((def_6_9<<1'd1) | ex_input0[14]) - (ex_input1[5:0] & {5'd6{jud_6_10}});
assign def_6_11 = ((def_6_10<<1'd1) | ex_input0[13]) - (ex_input1[5:0] & {5'd6{jud_6_11}});
assign def_6_12 = ((def_6_11<<1'd1) | ex_input0[12]) - (ex_input1[5:0] & {5'd6{jud_6_12}});
assign def_6_13 = ((def_6_12<<1'd1) | ex_input0[11]) - (ex_input1[5:0] & {5'd6{jud_6_13}});
assign def_6_14 = ((def_6_13<<1'd1) | ex_input0[10]) - (ex_input1[5:0] & {5'd6{jud_6_14}});
assign def_6_15 = ((def_6_14<<1'd1) | ex_input0[9]) - (ex_input1[5:0] & {5'd6{jud_6_15}});
assign def_6_16 = ((def_6_15<<1'd1) | ex_input0[8]) - (ex_input1[5:0] & {5'd6{jud_6_16}});
assign def_6_17 = ((def_6_16<<1'd1) | ex_input0[7]) - (ex_input1[5:0] & {5'd6{jud_6_17}});
assign def_6_18 = ((def_6_17<<1'd1) | ex_input0[6]) - (ex_input1[5:0] & {5'd6{jud_6_18}});
assign def_6_19 = ((def_6_18<<1'd1) | ex_input0[5]) - (ex_input1[5:0] & {5'd6{jud_6_19}});
assign def_6_20 = ((def_6_19<<1'd1) | ex_input0[4]) - (ex_input1[5:0] & {5'd6{jud_6_20}});
assign def_6_21 = ((def_6_20<<1'd1) | ex_input0[3]) - (ex_input1[5:0] & {5'd6{jud_6_21}});
assign def_6_22 = ((def_6_21<<1'd1) | ex_input0[2]) - (ex_input1[5:0] & {5'd6{jud_6_22}});
assign def_6_23 = ((def_6_22<<1'd1) | ex_input0[1]) - (ex_input1[5:0] & {5'd6{jud_6_23}});
assign def_6_24 = ((def_6_23<<1'd1) | ex_input0[0]) - (ex_input1[5:0] & {5'd6{jud_6_24}});

assign ans_6[29] = 1'd0;
assign ans_6[28] = 1'd0;
assign ans_6[27] = 1'd0;
assign ans_6[26] = 1'd0;
assign ans_6[25] = 1'd0;
assign ans_6[24] = jud_6_0;
assign ans_6[23] = jud_6_1;
assign ans_6[22] = jud_6_2;
assign ans_6[21] = jud_6_3;
assign ans_6[20] = jud_6_4;
assign ans_6[19] = jud_6_5;
assign ans_6[18] = jud_6_6;
assign ans_6[17] = jud_6_7;
assign ans_6[16] = jud_6_8;
assign ans_6[15] = jud_6_9;
assign ans_6[14] = jud_6_10;
assign ans_6[13] = jud_6_11;
assign ans_6[12] = jud_6_12;
assign ans_6[11] = jud_6_13;
assign ans_6[10] = jud_6_14;
assign ans_6[9] = jud_6_15;
assign ans_6[8] = jud_6_16;
assign ans_6[7] = jud_6_17;
assign ans_6[6] = jud_6_18;
assign ans_6[5] = jud_6_19;
assign ans_6[4] = jud_6_20;
assign ans_6[3] = jud_6_21;
assign ans_6[2] = jud_6_22;
assign ans_6[1] = jud_6_23;
assign ans_6[0] = jud_6_24;

//  5bit /////////////////////////////////////////////////////////////////////////////
assign jud_5_0 = ex_input0[29:25] >= ex_input1[4:0];
assign jud_5_1 = ((def_5_0<<1'd1) | ex_input0[24]) >= ex_input1[4:0];
assign jud_5_2 = ((def_5_1<<1'd1) | ex_input0[23]) >= ex_input1[4:0];
assign jud_5_3 = ((def_5_2<<1'd1) | ex_input0[22]) >= ex_input1[4:0];
assign jud_5_4 = ((def_5_3<<1'd1) | ex_input0[21]) >= ex_input1[4:0];
assign jud_5_5 = ((def_5_4<<1'd1) | ex_input0[20]) >= ex_input1[4:0];
assign jud_5_6 = ((def_5_5<<1'd1) | ex_input0[19]) >= ex_input1[4:0];
assign jud_5_7 = ((def_5_6<<1'd1) | ex_input0[18]) >= ex_input1[4:0];
assign jud_5_8 = ((def_5_7<<1'd1) | ex_input0[17]) >= ex_input1[4:0];
assign jud_5_9 = ((def_5_8<<1'd1) | ex_input0[16]) >= ex_input1[4:0];
assign jud_5_10 = ((def_5_9<<1'd1) | ex_input0[15]) >= ex_input1[4:0];
assign jud_5_11 = ((def_5_10<<1'd1) | ex_input0[14]) >= ex_input1[4:0];
assign jud_5_12 = ((def_5_11<<1'd1) | ex_input0[13]) >= ex_input1[4:0];
assign jud_5_13 = ((def_5_12<<1'd1) | ex_input0[12]) >= ex_input1[4:0];
assign jud_5_14 = ((def_5_13<<1'd1) | ex_input0[11]) >= ex_input1[4:0];
assign jud_5_15 = ((def_5_14<<1'd1) | ex_input0[10]) >= ex_input1[4:0];
assign jud_5_16 = ((def_5_15<<1'd1) | ex_input0[9]) >= ex_input1[4:0];
assign jud_5_17 = ((def_5_16<<1'd1) | ex_input0[8]) >= ex_input1[4:0];
assign jud_5_18 = ((def_5_17<<1'd1) | ex_input0[7]) >= ex_input1[4:0];
assign jud_5_19 = ((def_5_18<<1'd1) | ex_input0[6]) >= ex_input1[4:0];
assign jud_5_20 = ((def_5_19<<1'd1) | ex_input0[5]) >= ex_input1[4:0];
assign jud_5_21 = ((def_5_20<<1'd1) | ex_input0[4]) >= ex_input1[4:0];
assign jud_5_22 = ((def_5_21<<1'd1) | ex_input0[3]) >= ex_input1[4:0];
assign jud_5_23 = ((def_5_22<<1'd1) | ex_input0[2]) >= ex_input1[4:0];
assign jud_5_24 = ((def_5_23<<1'd1) | ex_input0[1]) >= ex_input1[4:0];
assign jud_5_25 = ((def_5_24<<1'd1) | ex_input0[0]) >= ex_input1[4:0];

assign def_5_0 = ex_input0[29:25] - (ex_input1[4:0] & {5'd5{jud_5_0}});
assign def_5_1 = ((def_5_0<<1'd1) | ex_input0[24]) - (ex_input1[4:0] & {5'd5{jud_5_1}});
assign def_5_2 = ((def_5_1<<1'd1) | ex_input0[23]) - (ex_input1[4:0] & {5'd5{jud_5_2}});
assign def_5_3 = ((def_5_2<<1'd1) | ex_input0[22]) - (ex_input1[4:0] & {5'd5{jud_5_3}});
assign def_5_4 = ((def_5_3<<1'd1) | ex_input0[21]) - (ex_input1[4:0] & {5'd5{jud_5_4}});
assign def_5_5 = ((def_5_4<<1'd1) | ex_input0[20]) - (ex_input1[4:0] & {5'd5{jud_5_5}});
assign def_5_6 = ((def_5_5<<1'd1) | ex_input0[19]) - (ex_input1[4:0] & {5'd5{jud_5_6}});
assign def_5_7 = ((def_5_6<<1'd1) | ex_input0[18]) - (ex_input1[4:0] & {5'd5{jud_5_7}});
assign def_5_8 = ((def_5_7<<1'd1) | ex_input0[17]) - (ex_input1[4:0] & {5'd5{jud_5_8}});
assign def_5_9 = ((def_5_8<<1'd1) | ex_input0[16]) - (ex_input1[4:0] & {5'd5{jud_5_9}});
assign def_5_10 = ((def_5_9<<1'd1) | ex_input0[15]) - (ex_input1[4:0] & {5'd5{jud_5_10}});
assign def_5_11 = ((def_5_10<<1'd1) | ex_input0[14]) - (ex_input1[4:0] & {5'd5{jud_5_11}});
assign def_5_12 = ((def_5_11<<1'd1) | ex_input0[13]) - (ex_input1[4:0] & {5'd5{jud_5_12}});
assign def_5_13 = ((def_5_12<<1'd1) | ex_input0[12]) - (ex_input1[4:0] & {5'd5{jud_5_13}});
assign def_5_14 = ((def_5_13<<1'd1) | ex_input0[11]) - (ex_input1[4:0] & {5'd5{jud_5_14}});
assign def_5_15 = ((def_5_14<<1'd1) | ex_input0[10]) - (ex_input1[4:0] & {5'd5{jud_5_15}});
assign def_5_16 = ((def_5_15<<1'd1) | ex_input0[9]) - (ex_input1[4:0] & {5'd5{jud_5_16}});
assign def_5_17 = ((def_5_16<<1'd1) | ex_input0[8]) - (ex_input1[4:0] & {5'd5{jud_5_17}});
assign def_5_18 = ((def_5_17<<1'd1) | ex_input0[7]) - (ex_input1[4:0] & {5'd5{jud_5_18}});
assign def_5_19 = ((def_5_18<<1'd1) | ex_input0[6]) - (ex_input1[4:0] & {5'd5{jud_5_19}});
assign def_5_20 = ((def_5_19<<1'd1) | ex_input0[5]) - (ex_input1[4:0] & {5'd5{jud_5_20}});
assign def_5_21 = ((def_5_20<<1'd1) | ex_input0[4]) - (ex_input1[4:0] & {5'd5{jud_5_21}});
assign def_5_22 = ((def_5_21<<1'd1) | ex_input0[3]) - (ex_input1[4:0] & {5'd5{jud_5_22}});
assign def_5_23 = ((def_5_22<<1'd1) | ex_input0[2]) - (ex_input1[4:0] & {5'd5{jud_5_23}});
assign def_5_24 = ((def_5_23<<1'd1) | ex_input0[1]) - (ex_input1[4:0] & {5'd5{jud_5_24}});
assign def_5_25 = ((def_5_24<<1'd1) | ex_input0[0]) - (ex_input1[4:0] & {5'd5{jud_5_25}});

assign ans_5[29] = 1'd0;
assign ans_5[28] = 1'd0;
assign ans_5[27] = 1'd0;
assign ans_5[26] = 1'd0;
assign ans_5[25] = jud_5_0;
assign ans_5[24] = jud_5_1;
assign ans_5[23] = jud_5_2;
assign ans_5[22] = jud_5_3;
assign ans_5[21] = jud_5_4;
assign ans_5[20] = jud_5_5;
assign ans_5[19] = jud_5_6;
assign ans_5[18] = jud_5_7;
assign ans_5[17] = jud_5_8;
assign ans_5[16] = jud_5_9;
assign ans_5[15] = jud_5_10;
assign ans_5[14] = jud_5_11;
assign ans_5[13] = jud_5_12;
assign ans_5[12] = jud_5_13;
assign ans_5[11] = jud_5_14;
assign ans_5[10] = jud_5_15;
assign ans_5[9] = jud_5_16;
assign ans_5[8] = jud_5_17;
assign ans_5[7] = jud_5_18;
assign ans_5[6] = jud_5_19;
assign ans_5[5] = jud_5_20;
assign ans_5[4] = jud_5_21;
assign ans_5[3] = jud_5_22;
assign ans_5[2] = jud_5_23;
assign ans_5[1] = jud_5_24;
assign ans_5[0] = jud_5_25;

//  4bit /////////////////////////////////////////////////////////////////////////////
assign jud_4_0 = ex_input0[29:26] >= ex_input1[3:0];
assign jud_4_1 = ((def_4_0<<1'd1) | ex_input0[25]) >= ex_input1[3:0];
assign jud_4_2 = ((def_4_1<<1'd1) | ex_input0[24]) >= ex_input1[3:0];
assign jud_4_3 = ((def_4_2<<1'd1) | ex_input0[23]) >= ex_input1[3:0];
assign jud_4_4 = ((def_4_3<<1'd1) | ex_input0[22]) >= ex_input1[3:0];
assign jud_4_5 = ((def_4_4<<1'd1) | ex_input0[21]) >= ex_input1[3:0];
assign jud_4_6 = ((def_4_5<<1'd1) | ex_input0[20]) >= ex_input1[3:0];
assign jud_4_7 = ((def_4_6<<1'd1) | ex_input0[19]) >= ex_input1[3:0];
assign jud_4_8 = ((def_4_7<<1'd1) | ex_input0[18]) >= ex_input1[3:0];
assign jud_4_9 = ((def_4_8<<1'd1) | ex_input0[17]) >= ex_input1[3:0];
assign jud_4_10 = ((def_4_9<<1'd1) | ex_input0[16]) >= ex_input1[3:0];
assign jud_4_11 = ((def_4_10<<1'd1) | ex_input0[15]) >= ex_input1[3:0];
assign jud_4_12 = ((def_4_11<<1'd1) | ex_input0[14]) >= ex_input1[3:0];
assign jud_4_13 = ((def_4_12<<1'd1) | ex_input0[13]) >= ex_input1[3:0];
assign jud_4_14 = ((def_4_13<<1'd1) | ex_input0[12]) >= ex_input1[3:0];
assign jud_4_15 = ((def_4_14<<1'd1) | ex_input0[11]) >= ex_input1[3:0];
assign jud_4_16 = ((def_4_15<<1'd1) | ex_input0[10]) >= ex_input1[3:0];
assign jud_4_17 = ((def_4_16<<1'd1) | ex_input0[9]) >= ex_input1[3:0];
assign jud_4_18 = ((def_4_17<<1'd1) | ex_input0[8]) >= ex_input1[3:0];
assign jud_4_19 = ((def_4_18<<1'd1) | ex_input0[7]) >= ex_input1[3:0];
assign jud_4_20 = ((def_4_19<<1'd1) | ex_input0[6]) >= ex_input1[3:0];
assign jud_4_21 = ((def_4_20<<1'd1) | ex_input0[5]) >= ex_input1[3:0];
assign jud_4_22 = ((def_4_21<<1'd1) | ex_input0[4]) >= ex_input1[3:0];
assign jud_4_23 = ((def_4_22<<1'd1) | ex_input0[3]) >= ex_input1[3:0];
assign jud_4_24 = ((def_4_23<<1'd1) | ex_input0[2]) >= ex_input1[3:0];
assign jud_4_25 = ((def_4_24<<1'd1) | ex_input0[1]) >= ex_input1[3:0];
assign jud_4_26 = ((def_4_25<<1'd1) | ex_input0[0]) >= ex_input1[3:0];

assign def_4_0 = ex_input0[29:26] - (ex_input1[3:0] & {5'd4{jud_4_0}});
assign def_4_1 = ((def_4_0<<1'd1) | ex_input0[25]) - (ex_input1[3:0] & {5'd4{jud_4_1}});
assign def_4_2 = ((def_4_1<<1'd1) | ex_input0[24]) - (ex_input1[3:0] & {5'd4{jud_4_2}});
assign def_4_3 = ((def_4_2<<1'd1) | ex_input0[23]) - (ex_input1[3:0] & {5'd4{jud_4_3}});
assign def_4_4 = ((def_4_3<<1'd1) | ex_input0[22]) - (ex_input1[3:0] & {5'd4{jud_4_4}});
assign def_4_5 = ((def_4_4<<1'd1) | ex_input0[21]) - (ex_input1[3:0] & {5'd4{jud_4_5}});
assign def_4_6 = ((def_4_5<<1'd1) | ex_input0[20]) - (ex_input1[3:0] & {5'd4{jud_4_6}});
assign def_4_7 = ((def_4_6<<1'd1) | ex_input0[19]) - (ex_input1[3:0] & {5'd4{jud_4_7}});
assign def_4_8 = ((def_4_7<<1'd1) | ex_input0[18]) - (ex_input1[3:0] & {5'd4{jud_4_8}});
assign def_4_9 = ((def_4_8<<1'd1) | ex_input0[17]) - (ex_input1[3:0] & {5'd4{jud_4_9}});
assign def_4_10 = ((def_4_9<<1'd1) | ex_input0[16]) - (ex_input1[3:0] & {5'd4{jud_4_10}});
assign def_4_11 = ((def_4_10<<1'd1) | ex_input0[15]) - (ex_input1[3:0] & {5'd4{jud_4_11}});
assign def_4_12 = ((def_4_11<<1'd1) | ex_input0[14]) - (ex_input1[3:0] & {5'd4{jud_4_12}});
assign def_4_13 = ((def_4_12<<1'd1) | ex_input0[13]) - (ex_input1[3:0] & {5'd4{jud_4_13}});
assign def_4_14 = ((def_4_13<<1'd1) | ex_input0[12]) - (ex_input1[3:0] & {5'd4{jud_4_14}});
assign def_4_15 = ((def_4_14<<1'd1) | ex_input0[11]) - (ex_input1[3:0] & {5'd4{jud_4_15}});
assign def_4_16 = ((def_4_15<<1'd1) | ex_input0[10]) - (ex_input1[3:0] & {5'd4{jud_4_16}});
assign def_4_17 = ((def_4_16<<1'd1) | ex_input0[9]) - (ex_input1[3:0] & {5'd4{jud_4_17}});
assign def_4_18 = ((def_4_17<<1'd1) | ex_input0[8]) - (ex_input1[3:0] & {5'd4{jud_4_18}});
assign def_4_19 = ((def_4_18<<1'd1) | ex_input0[7]) - (ex_input1[3:0] & {5'd4{jud_4_19}});
assign def_4_20 = ((def_4_19<<1'd1) | ex_input0[6]) - (ex_input1[3:0] & {5'd4{jud_4_20}});
assign def_4_21 = ((def_4_20<<1'd1) | ex_input0[5]) - (ex_input1[3:0] & {5'd4{jud_4_21}});
assign def_4_22 = ((def_4_21<<1'd1) | ex_input0[4]) - (ex_input1[3:0] & {5'd4{jud_4_22}});
assign def_4_23 = ((def_4_22<<1'd1) | ex_input0[3]) - (ex_input1[3:0] & {5'd4{jud_4_23}});
assign def_4_24 = ((def_4_23<<1'd1) | ex_input0[2]) - (ex_input1[3:0] & {5'd4{jud_4_24}});
assign def_4_25 = ((def_4_24<<1'd1) | ex_input0[1]) - (ex_input1[3:0] & {5'd4{jud_4_25}});
assign def_4_26 = ((def_4_25<<1'd1) | ex_input0[0]) - (ex_input1[3:0] & {5'd4{jud_4_26}});

assign ans_4[29] = 1'd0;
assign ans_4[28] = 1'd0;
assign ans_4[27] = 1'd0;
assign ans_4[26] = jud_4_0;
assign ans_4[25] = jud_4_1;
assign ans_4[24] = jud_4_2;
assign ans_4[23] = jud_4_3;
assign ans_4[22] = jud_4_4;
assign ans_4[21] = jud_4_5;
assign ans_4[20] = jud_4_6;
assign ans_4[19] = jud_4_7;
assign ans_4[18] = jud_4_8;
assign ans_4[17] = jud_4_9;
assign ans_4[16] = jud_4_10;
assign ans_4[15] = jud_4_11;
assign ans_4[14] = jud_4_12;
assign ans_4[13] = jud_4_13;
assign ans_4[12] = jud_4_14;
assign ans_4[11] = jud_4_15;
assign ans_4[10] = jud_4_16;
assign ans_4[9] = jud_4_17;
assign ans_4[8] = jud_4_18;
assign ans_4[7] = jud_4_19;
assign ans_4[6] = jud_4_20;
assign ans_4[5] = jud_4_21;
assign ans_4[4] = jud_4_22;
assign ans_4[3] = jud_4_23;
assign ans_4[2] = jud_4_24;
assign ans_4[1] = jud_4_25;
assign ans_4[0] = jud_4_26;

//  3bit /////////////////////////////////////////////////////////////////////////////
assign jud_3_0 = ex_input0[29:27] >= ex_input1[2:0];
assign jud_3_1 = ((def_3_0<<1'd1) | ex_input0[26]) >= ex_input1[2:0];
assign jud_3_2 = ((def_3_1<<1'd1) | ex_input0[25]) >= ex_input1[2:0];
assign jud_3_3 = ((def_3_2<<1'd1) | ex_input0[24]) >= ex_input1[2:0];
assign jud_3_4 = ((def_3_3<<1'd1) | ex_input0[23]) >= ex_input1[2:0];
assign jud_3_5 = ((def_3_4<<1'd1) | ex_input0[22]) >= ex_input1[2:0];
assign jud_3_6 = ((def_3_5<<1'd1) | ex_input0[21]) >= ex_input1[2:0];
assign jud_3_7 = ((def_3_6<<1'd1) | ex_input0[20]) >= ex_input1[2:0];
assign jud_3_8 = ((def_3_7<<1'd1) | ex_input0[19]) >= ex_input1[2:0];
assign jud_3_9 = ((def_3_8<<1'd1) | ex_input0[18]) >= ex_input1[2:0];
assign jud_3_10 = ((def_3_9<<1'd1) | ex_input0[17]) >= ex_input1[2:0];
assign jud_3_11 = ((def_3_10<<1'd1) | ex_input0[16]) >= ex_input1[2:0];
assign jud_3_12 = ((def_3_11<<1'd1) | ex_input0[15]) >= ex_input1[2:0];
assign jud_3_13 = ((def_3_12<<1'd1) | ex_input0[14]) >= ex_input1[2:0];
assign jud_3_14 = ((def_3_13<<1'd1) | ex_input0[13]) >= ex_input1[2:0];
assign jud_3_15 = ((def_3_14<<1'd1) | ex_input0[12]) >= ex_input1[2:0];
assign jud_3_16 = ((def_3_15<<1'd1) | ex_input0[11]) >= ex_input1[2:0];
assign jud_3_17 = ((def_3_16<<1'd1) | ex_input0[10]) >= ex_input1[2:0];
assign jud_3_18 = ((def_3_17<<1'd1) | ex_input0[9]) >= ex_input1[2:0];
assign jud_3_19 = ((def_3_18<<1'd1) | ex_input0[8]) >= ex_input1[2:0];
assign jud_3_20 = ((def_3_19<<1'd1) | ex_input0[7]) >= ex_input1[2:0];
assign jud_3_21 = ((def_3_20<<1'd1) | ex_input0[6]) >= ex_input1[2:0];
assign jud_3_22 = ((def_3_21<<1'd1) | ex_input0[5]) >= ex_input1[2:0];
assign jud_3_23 = ((def_3_22<<1'd1) | ex_input0[4]) >= ex_input1[2:0];
assign jud_3_24 = ((def_3_23<<1'd1) | ex_input0[3]) >= ex_input1[2:0];
assign jud_3_25 = ((def_3_24<<1'd1) | ex_input0[2]) >= ex_input1[2:0];
assign jud_3_26 = ((def_3_25<<1'd1) | ex_input0[1]) >= ex_input1[2:0];
assign jud_3_27 = ((def_3_26<<1'd1) | ex_input0[0]) >= ex_input1[2:0];

assign def_3_0 = ex_input0[29:27] - (ex_input1[2:0] & {5'd3{jud_3_0}});
assign def_3_1 = ((def_3_0<<1'd1) | ex_input0[26]) - (ex_input1[2:0] & {5'd3{jud_3_1}});
assign def_3_2 = ((def_3_1<<1'd1) | ex_input0[25]) - (ex_input1[2:0] & {5'd3{jud_3_2}});
assign def_3_3 = ((def_3_2<<1'd1) | ex_input0[24]) - (ex_input1[2:0] & {5'd3{jud_3_3}});
assign def_3_4 = ((def_3_3<<1'd1) | ex_input0[23]) - (ex_input1[2:0] & {5'd3{jud_3_4}});
assign def_3_5 = ((def_3_4<<1'd1) | ex_input0[22]) - (ex_input1[2:0] & {5'd3{jud_3_5}});
assign def_3_6 = ((def_3_5<<1'd1) | ex_input0[21]) - (ex_input1[2:0] & {5'd3{jud_3_6}});
assign def_3_7 = ((def_3_6<<1'd1) | ex_input0[20]) - (ex_input1[2:0] & {5'd3{jud_3_7}});
assign def_3_8 = ((def_3_7<<1'd1) | ex_input0[19]) - (ex_input1[2:0] & {5'd3{jud_3_8}});
assign def_3_9 = ((def_3_8<<1'd1) | ex_input0[18]) - (ex_input1[2:0] & {5'd3{jud_3_9}});
assign def_3_10 = ((def_3_9<<1'd1) | ex_input0[17]) - (ex_input1[2:0] & {5'd3{jud_3_10}});
assign def_3_11 = ((def_3_10<<1'd1) | ex_input0[16]) - (ex_input1[2:0] & {5'd3{jud_3_11}});
assign def_3_12 = ((def_3_11<<1'd1) | ex_input0[15]) - (ex_input1[2:0] & {5'd3{jud_3_12}});
assign def_3_13 = ((def_3_12<<1'd1) | ex_input0[14]) - (ex_input1[2:0] & {5'd3{jud_3_13}});
assign def_3_14 = ((def_3_13<<1'd1) | ex_input0[13]) - (ex_input1[2:0] & {5'd3{jud_3_14}});
assign def_3_15 = ((def_3_14<<1'd1) | ex_input0[12]) - (ex_input1[2:0] & {5'd3{jud_3_15}});
assign def_3_16 = ((def_3_15<<1'd1) | ex_input0[11]) - (ex_input1[2:0] & {5'd3{jud_3_16}});
assign def_3_17 = ((def_3_16<<1'd1) | ex_input0[10]) - (ex_input1[2:0] & {5'd3{jud_3_17}});
assign def_3_18 = ((def_3_17<<1'd1) | ex_input0[9]) - (ex_input1[2:0] & {5'd3{jud_3_18}});
assign def_3_19 = ((def_3_18<<1'd1) | ex_input0[8]) - (ex_input1[2:0] & {5'd3{jud_3_19}});
assign def_3_20 = ((def_3_19<<1'd1) | ex_input0[7]) - (ex_input1[2:0] & {5'd3{jud_3_20}});
assign def_3_21 = ((def_3_20<<1'd1) | ex_input0[6]) - (ex_input1[2:0] & {5'd3{jud_3_21}});
assign def_3_22 = ((def_3_21<<1'd1) | ex_input0[5]) - (ex_input1[2:0] & {5'd3{jud_3_22}});
assign def_3_23 = ((def_3_22<<1'd1) | ex_input0[4]) - (ex_input1[2:0] & {5'd3{jud_3_23}});
assign def_3_24 = ((def_3_23<<1'd1) | ex_input0[3]) - (ex_input1[2:0] & {5'd3{jud_3_24}});
assign def_3_25 = ((def_3_24<<1'd1) | ex_input0[2]) - (ex_input1[2:0] & {5'd3{jud_3_25}});
assign def_3_26 = ((def_3_25<<1'd1) | ex_input0[1]) - (ex_input1[2:0] & {5'd3{jud_3_26}});
assign def_3_27 = ((def_3_26<<1'd1) | ex_input0[0]) - (ex_input1[2:0] & {5'd3{jud_3_27}});

assign ans_3[29] = 1'd0;
assign ans_3[28] = 1'd0;
assign ans_3[27] = jud_3_0;
assign ans_3[26] = jud_3_1;
assign ans_3[25] = jud_3_2;
assign ans_3[24] = jud_3_3;
assign ans_3[23] = jud_3_4;
assign ans_3[22] = jud_3_5;
assign ans_3[21] = jud_3_6;
assign ans_3[20] = jud_3_7;
assign ans_3[19] = jud_3_8;
assign ans_3[18] = jud_3_9;
assign ans_3[17] = jud_3_10;
assign ans_3[16] = jud_3_11;
assign ans_3[15] = jud_3_12;
assign ans_3[14] = jud_3_13;
assign ans_3[13] = jud_3_14;
assign ans_3[12] = jud_3_15;
assign ans_3[11] = jud_3_16;
assign ans_3[10] = jud_3_17;
assign ans_3[9] = jud_3_18;
assign ans_3[8] = jud_3_19;
assign ans_3[7] = jud_3_20;
assign ans_3[6] = jud_3_21;
assign ans_3[5] = jud_3_22;
assign ans_3[4] = jud_3_23;
assign ans_3[3] = jud_3_24;
assign ans_3[2] = jud_3_25;
assign ans_3[1] = jud_3_26;
assign ans_3[0] = jud_3_27;

//  2bit /////////////////////////////////////////////////////////////////////////////
assign jud_2_0 = ex_input0[29:28] >= ex_input1[1:0];
assign jud_2_1 = ((def_2_0<<1'd1) | ex_input0[27]) >= ex_input1[1:0];
assign jud_2_2 = ((def_2_1<<1'd1) | ex_input0[26]) >= ex_input1[1:0];
assign jud_2_3 = ((def_2_2<<1'd1) | ex_input0[25]) >= ex_input1[1:0];
assign jud_2_4 = ((def_2_3<<1'd1) | ex_input0[24]) >= ex_input1[1:0];
assign jud_2_5 = ((def_2_4<<1'd1) | ex_input0[23]) >= ex_input1[1:0];
assign jud_2_6 = ((def_2_5<<1'd1) | ex_input0[22]) >= ex_input1[1:0];
assign jud_2_7 = ((def_2_6<<1'd1) | ex_input0[21]) >= ex_input1[1:0];
assign jud_2_8 = ((def_2_7<<1'd1) | ex_input0[20]) >= ex_input1[1:0];
assign jud_2_9 = ((def_2_8<<1'd1) | ex_input0[19]) >= ex_input1[1:0];
assign jud_2_10 = ((def_2_9<<1'd1) | ex_input0[18]) >= ex_input1[1:0];
assign jud_2_11 = ((def_2_10<<1'd1) | ex_input0[17]) >= ex_input1[1:0];
assign jud_2_12 = ((def_2_11<<1'd1) | ex_input0[16]) >= ex_input1[1:0];
assign jud_2_13 = ((def_2_12<<1'd1) | ex_input0[15]) >= ex_input1[1:0];
assign jud_2_14 = ((def_2_13<<1'd1) | ex_input0[14]) >= ex_input1[1:0];
assign jud_2_15 = ((def_2_14<<1'd1) | ex_input0[13]) >= ex_input1[1:0];
assign jud_2_16 = ((def_2_15<<1'd1) | ex_input0[12]) >= ex_input1[1:0];
assign jud_2_17 = ((def_2_16<<1'd1) | ex_input0[11]) >= ex_input1[1:0];
assign jud_2_18 = ((def_2_17<<1'd1) | ex_input0[10]) >= ex_input1[1:0];
assign jud_2_19 = ((def_2_18<<1'd1) | ex_input0[9]) >= ex_input1[1:0];
assign jud_2_20 = ((def_2_19<<1'd1) | ex_input0[8]) >= ex_input1[1:0];
assign jud_2_21 = ((def_2_20<<1'd1) | ex_input0[7]) >= ex_input1[1:0];
assign jud_2_22 = ((def_2_21<<1'd1) | ex_input0[6]) >= ex_input1[1:0];
assign jud_2_23 = ((def_2_22<<1'd1) | ex_input0[5]) >= ex_input1[1:0];
assign jud_2_24 = ((def_2_23<<1'd1) | ex_input0[4]) >= ex_input1[1:0];
assign jud_2_25 = ((def_2_24<<1'd1) | ex_input0[3]) >= ex_input1[1:0];
assign jud_2_26 = ((def_2_25<<1'd1) | ex_input0[2]) >= ex_input1[1:0];
assign jud_2_27 = ((def_2_26<<1'd1) | ex_input0[1]) >= ex_input1[1:0];
assign jud_2_28 = ((def_2_27<<1'd1) | ex_input0[0]) >= ex_input1[1:0];

assign def_2_0 = ex_input0[29:28] - (ex_input1[1:0] & {5'd2{jud_2_0}});
assign def_2_1 = ((def_2_0<<1'd1) | ex_input0[27]) - (ex_input1[1:0] & {5'd2{jud_2_1}});
assign def_2_2 = ((def_2_1<<1'd1) | ex_input0[26]) - (ex_input1[1:0] & {5'd2{jud_2_2}});
assign def_2_3 = ((def_2_2<<1'd1) | ex_input0[25]) - (ex_input1[1:0] & {5'd2{jud_2_3}});
assign def_2_4 = ((def_2_3<<1'd1) | ex_input0[24]) - (ex_input1[1:0] & {5'd2{jud_2_4}});
assign def_2_5 = ((def_2_4<<1'd1) | ex_input0[23]) - (ex_input1[1:0] & {5'd2{jud_2_5}});
assign def_2_6 = ((def_2_5<<1'd1) | ex_input0[22]) - (ex_input1[1:0] & {5'd2{jud_2_6}});
assign def_2_7 = ((def_2_6<<1'd1) | ex_input0[21]) - (ex_input1[1:0] & {5'd2{jud_2_7}});
assign def_2_8 = ((def_2_7<<1'd1) | ex_input0[20]) - (ex_input1[1:0] & {5'd2{jud_2_8}});
assign def_2_9 = ((def_2_8<<1'd1) | ex_input0[19]) - (ex_input1[1:0] & {5'd2{jud_2_9}});
assign def_2_10 = ((def_2_9<<1'd1) | ex_input0[18]) - (ex_input1[1:0] & {5'd2{jud_2_10}});
assign def_2_11 = ((def_2_10<<1'd1) | ex_input0[17]) - (ex_input1[1:0] & {5'd2{jud_2_11}});
assign def_2_12 = ((def_2_11<<1'd1) | ex_input0[16]) - (ex_input1[1:0] & {5'd2{jud_2_12}});
assign def_2_13 = ((def_2_12<<1'd1) | ex_input0[15]) - (ex_input1[1:0] & {5'd2{jud_2_13}});
assign def_2_14 = ((def_2_13<<1'd1) | ex_input0[14]) - (ex_input1[1:0] & {5'd2{jud_2_14}});
assign def_2_15 = ((def_2_14<<1'd1) | ex_input0[13]) - (ex_input1[1:0] & {5'd2{jud_2_15}});
assign def_2_16 = ((def_2_15<<1'd1) | ex_input0[12]) - (ex_input1[1:0] & {5'd2{jud_2_16}});
assign def_2_17 = ((def_2_16<<1'd1) | ex_input0[11]) - (ex_input1[1:0] & {5'd2{jud_2_17}});
assign def_2_18 = ((def_2_17<<1'd1) | ex_input0[10]) - (ex_input1[1:0] & {5'd2{jud_2_18}});
assign def_2_19 = ((def_2_18<<1'd1) | ex_input0[9]) - (ex_input1[1:0] & {5'd2{jud_2_19}});
assign def_2_20 = ((def_2_19<<1'd1) | ex_input0[8]) - (ex_input1[1:0] & {5'd2{jud_2_20}});
assign def_2_21 = ((def_2_20<<1'd1) | ex_input0[7]) - (ex_input1[1:0] & {5'd2{jud_2_21}});
assign def_2_22 = ((def_2_21<<1'd1) | ex_input0[6]) - (ex_input1[1:0] & {5'd2{jud_2_22}});
assign def_2_23 = ((def_2_22<<1'd1) | ex_input0[5]) - (ex_input1[1:0] & {5'd2{jud_2_23}});
assign def_2_24 = ((def_2_23<<1'd1) | ex_input0[4]) - (ex_input1[1:0] & {5'd2{jud_2_24}});
assign def_2_25 = ((def_2_24<<1'd1) | ex_input0[3]) - (ex_input1[1:0] & {5'd2{jud_2_25}});
assign def_2_26 = ((def_2_25<<1'd1) | ex_input0[2]) - (ex_input1[1:0] & {5'd2{jud_2_26}});
assign def_2_27 = ((def_2_26<<1'd1) | ex_input0[1]) - (ex_input1[1:0] & {5'd2{jud_2_27}});
assign def_2_28 = ((def_2_27<<1'd1) | ex_input0[0]) - (ex_input1[1:0] & {5'd2{jud_2_28}});

assign ans_2[29] = 1'd0;
assign ans_2[28] = jud_2_0;
assign ans_2[27] = jud_2_1;
assign ans_2[26] = jud_2_2;
assign ans_2[25] = jud_2_3;
assign ans_2[24] = jud_2_4;
assign ans_2[23] = jud_2_5;
assign ans_2[22] = jud_2_6;
assign ans_2[21] = jud_2_7;
assign ans_2[20] = jud_2_8;
assign ans_2[19] = jud_2_9;
assign ans_2[18] = jud_2_10;
assign ans_2[17] = jud_2_11;
assign ans_2[16] = jud_2_12;
assign ans_2[15] = jud_2_13;
assign ans_2[14] = jud_2_14;
assign ans_2[13] = jud_2_15;
assign ans_2[12] = jud_2_16;
assign ans_2[11] = jud_2_17;
assign ans_2[10] = jud_2_18;
assign ans_2[9] = jud_2_19;
assign ans_2[8] = jud_2_20;
assign ans_2[7] = jud_2_21;
assign ans_2[6] = jud_2_22;
assign ans_2[5] = jud_2_23;
assign ans_2[4] = jud_2_24;
assign ans_2[3] = jud_2_25;
assign ans_2[2] = jud_2_26;
assign ans_2[1] = jud_2_27;
assign ans_2[0] = jud_2_28;

//  1bit /////////////////////////////////////////////////////////////////////////////
assign jud_1_0 = ex_input0[29] >= ex_input1[0];
assign jud_1_1 = ((def_1_0<<1'd1) | ex_input0[28]) >= ex_input1[0];
assign jud_1_2 = ((def_1_1<<1'd1) | ex_input0[27]) >= ex_input1[0];
assign jud_1_3 = ((def_1_2<<1'd1) | ex_input0[26]) >= ex_input1[0];
assign jud_1_4 = ((def_1_3<<1'd1) | ex_input0[25]) >= ex_input1[0];
assign jud_1_5 = ((def_1_4<<1'd1) | ex_input0[24]) >= ex_input1[0];
assign jud_1_6 = ((def_1_5<<1'd1) | ex_input0[23]) >= ex_input1[0];
assign jud_1_7 = ((def_1_6<<1'd1) | ex_input0[22]) >= ex_input1[0];
assign jud_1_8 = ((def_1_7<<1'd1) | ex_input0[21]) >= ex_input1[0];
assign jud_1_9 = ((def_1_8<<1'd1) | ex_input0[20]) >= ex_input1[0];
assign jud_1_10 = ((def_1_9<<1'd1) | ex_input0[19]) >= ex_input1[0];
assign jud_1_11 = ((def_1_10<<1'd1) | ex_input0[18]) >= ex_input1[0];
assign jud_1_12 = ((def_1_11<<1'd1) | ex_input0[17]) >= ex_input1[0];
assign jud_1_13 = ((def_1_12<<1'd1) | ex_input0[16]) >= ex_input1[0];
assign jud_1_14 = ((def_1_13<<1'd1) | ex_input0[15]) >= ex_input1[0];
assign jud_1_15 = ((def_1_14<<1'd1) | ex_input0[14]) >= ex_input1[0];
assign jud_1_16 = ((def_1_15<<1'd1) | ex_input0[13]) >= ex_input1[0];
assign jud_1_17 = ((def_1_16<<1'd1) | ex_input0[12]) >= ex_input1[0];
assign jud_1_18 = ((def_1_17<<1'd1) | ex_input0[11]) >= ex_input1[0];
assign jud_1_19 = ((def_1_18<<1'd1) | ex_input0[10]) >= ex_input1[0];
assign jud_1_20 = ((def_1_19<<1'd1) | ex_input0[9]) >= ex_input1[0];
assign jud_1_21 = ((def_1_20<<1'd1) | ex_input0[8]) >= ex_input1[0];
assign jud_1_22 = ((def_1_21<<1'd1) | ex_input0[7]) >= ex_input1[0];
assign jud_1_23 = ((def_1_22<<1'd1) | ex_input0[6]) >= ex_input1[0];
assign jud_1_24 = ((def_1_23<<1'd1) | ex_input0[5]) >= ex_input1[0];
assign jud_1_25 = ((def_1_24<<1'd1) | ex_input0[4]) >= ex_input1[0];
assign jud_1_26 = ((def_1_25<<1'd1) | ex_input0[3]) >= ex_input1[0];
assign jud_1_27 = ((def_1_26<<1'd1) | ex_input0[2]) >= ex_input1[0];
assign jud_1_28 = ((def_1_27<<1'd1) | ex_input0[1]) >= ex_input1[0];
assign jud_1_29 = ((def_1_28<<1'd1) | ex_input0[0]) >= ex_input1[0];

assign def_1_0 = ex_input0[29] - (ex_input1[0] & {5'd1{jud_1_0}});
assign def_1_1 = ((def_1_0<<1'd1) | ex_input0[28]) - (ex_input1[0] & {5'd1{jud_1_1}});
assign def_1_2 = ((def_1_1<<1'd1) | ex_input0[27]) - (ex_input1[0] & {5'd1{jud_1_2}});
assign def_1_3 = ((def_1_2<<1'd1) | ex_input0[26]) - (ex_input1[0] & {5'd1{jud_1_3}});
assign def_1_4 = ((def_1_3<<1'd1) | ex_input0[25]) - (ex_input1[0] & {5'd1{jud_1_4}});
assign def_1_5 = ((def_1_4<<1'd1) | ex_input0[24]) - (ex_input1[0] & {5'd1{jud_1_5}});
assign def_1_6 = ((def_1_5<<1'd1) | ex_input0[23]) - (ex_input1[0] & {5'd1{jud_1_6}});
assign def_1_7 = ((def_1_6<<1'd1) | ex_input0[22]) - (ex_input1[0] & {5'd1{jud_1_7}});
assign def_1_8 = ((def_1_7<<1'd1) | ex_input0[21]) - (ex_input1[0] & {5'd1{jud_1_8}});
assign def_1_9 = ((def_1_8<<1'd1) | ex_input0[20]) - (ex_input1[0] & {5'd1{jud_1_9}});
assign def_1_10 = ((def_1_9<<1'd1) | ex_input0[19]) - (ex_input1[0] & {5'd1{jud_1_10}});
assign def_1_11 = ((def_1_10<<1'd1) | ex_input0[18]) - (ex_input1[0] & {5'd1{jud_1_11}});
assign def_1_12 = ((def_1_11<<1'd1) | ex_input0[17]) - (ex_input1[0] & {5'd1{jud_1_12}});
assign def_1_13 = ((def_1_12<<1'd1) | ex_input0[16]) - (ex_input1[0] & {5'd1{jud_1_13}});
assign def_1_14 = ((def_1_13<<1'd1) | ex_input0[15]) - (ex_input1[0] & {5'd1{jud_1_14}});
assign def_1_15 = ((def_1_14<<1'd1) | ex_input0[14]) - (ex_input1[0] & {5'd1{jud_1_15}});
assign def_1_16 = ((def_1_15<<1'd1) | ex_input0[13]) - (ex_input1[0] & {5'd1{jud_1_16}});
assign def_1_17 = ((def_1_16<<1'd1) | ex_input0[12]) - (ex_input1[0] & {5'd1{jud_1_17}});
assign def_1_18 = ((def_1_17<<1'd1) | ex_input0[11]) - (ex_input1[0] & {5'd1{jud_1_18}});
assign def_1_19 = ((def_1_18<<1'd1) | ex_input0[10]) - (ex_input1[0] & {5'd1{jud_1_19}});
assign def_1_20 = ((def_1_19<<1'd1) | ex_input0[9]) - (ex_input1[0] & {5'd1{jud_1_20}});
assign def_1_21 = ((def_1_20<<1'd1) | ex_input0[8]) - (ex_input1[0] & {5'd1{jud_1_21}});
assign def_1_22 = ((def_1_21<<1'd1) | ex_input0[7]) - (ex_input1[0] & {5'd1{jud_1_22}});
assign def_1_23 = ((def_1_22<<1'd1) | ex_input0[6]) - (ex_input1[0] & {5'd1{jud_1_23}});
assign def_1_24 = ((def_1_23<<1'd1) | ex_input0[5]) - (ex_input1[0] & {5'd1{jud_1_24}});
assign def_1_25 = ((def_1_24<<1'd1) | ex_input0[4]) - (ex_input1[0] & {5'd1{jud_1_25}});
assign def_1_26 = ((def_1_25<<1'd1) | ex_input0[3]) - (ex_input1[0] & {5'd1{jud_1_26}});
assign def_1_27 = ((def_1_26<<1'd1) | ex_input0[2]) - (ex_input1[0] & {5'd1{jud_1_27}});
assign def_1_28 = ((def_1_27<<1'd1) | ex_input0[1]) - (ex_input1[0] & {5'd1{jud_1_28}});
assign def_1_29 = ((def_1_28<<1'd1) | ex_input0[0]) - (ex_input1[0] & {5'd1{jud_1_29}});

assign ans_1[29] = jud_1_0;
assign ans_1[28] = jud_1_1;
assign ans_1[27] = jud_1_2;
assign ans_1[26] = jud_1_3;
assign ans_1[25] = jud_1_4;
assign ans_1[24] = jud_1_5;
assign ans_1[23] = jud_1_6;
assign ans_1[22] = jud_1_7;
assign ans_1[21] = jud_1_8;
assign ans_1[20] = jud_1_9;
assign ans_1[19] = jud_1_10;
assign ans_1[18] = jud_1_11;
assign ans_1[17] = jud_1_12;
assign ans_1[16] = jud_1_13;
assign ans_1[15] = jud_1_14;
assign ans_1[14] = jud_1_15;
assign ans_1[13] = jud_1_16;
assign ans_1[12] = jud_1_17;
assign ans_1[11] = jud_1_18;
assign ans_1[10] = jud_1_19;
assign ans_1[9] = jud_1_20;
assign ans_1[8] = jud_1_21;
assign ans_1[7] = jud_1_22;
assign ans_1[6] = jud_1_23;
assign ans_1[5] = jud_1_24;
assign ans_1[4] = jud_1_25;
assign ans_1[3] = jud_1_26;
assign ans_1[2] = jud_1_27;
assign ans_1[1] = jud_1_28;
assign ans_1[0] = jud_1_29;



assign msb_20 = (INPUT_1[19]&(~INPUT_0[20])) | (comp_input1[19]&INPUT_0[20]);
assign msb_19 = (INPUT_1[18]&(~INPUT_0[20])) | (comp_input1[18]&INPUT_0[20]);
assign msb_18 = (INPUT_1[17]&(~INPUT_0[20])) | (comp_input1[17]&INPUT_0[20]);
assign msb_17 = (INPUT_1[16]&(~INPUT_0[20])) | (comp_input1[16]&INPUT_0[20]);
assign msb_16 = (INPUT_1[15]&(~INPUT_0[20])) | (comp_input1[15]&INPUT_0[20]);
assign msb_15 = (INPUT_1[14]&(~INPUT_0[20])) | (comp_input1[14]&INPUT_0[20]);
assign msb_14 = (INPUT_1[13]&(~INPUT_0[20])) | (comp_input1[13]&INPUT_0[20]);
assign msb_13 = (INPUT_1[12]&(~INPUT_0[20])) | (comp_input1[12]&INPUT_0[20]);
assign msb_12 = (INPUT_1[11]&(~INPUT_0[20])) | (comp_input1[11]&INPUT_0[20]);
assign msb_11 = (INPUT_1[10]&(~INPUT_0[20])) | (comp_input1[10]&INPUT_0[20]);
assign msb_10 = (INPUT_1[9]&(~INPUT_0[20])) | (comp_input1[9]&INPUT_0[20]);
assign msb_9 = (INPUT_1[8]&(~INPUT_0[20])) | (comp_input1[8]&INPUT_0[20]);
assign msb_8 = (INPUT_1[7]&(~INPUT_0[20])) | (comp_input1[7]&INPUT_0[20]);
assign msb_7 = (INPUT_1[6]&(~INPUT_0[20])) | (comp_input1[6]&INPUT_0[20]);
assign msb_6 = (INPUT_1[5]&(~INPUT_0[20])) | (comp_input1[5]&INPUT_0[20]);
assign msb_5 = (INPUT_1[4]&(~INPUT_0[20])) | (comp_input1[4]&INPUT_0[20]);
assign msb_4 = (INPUT_1[3]&(~INPUT_0[20])) | (comp_input1[3]&INPUT_0[20]);
assign msb_3 = (INPUT_1[2]&(~INPUT_0[20])) | (comp_input1[2]&INPUT_0[20]);
assign msb_2 = (INPUT_1[1]&(~INPUT_0[20])) | (comp_input1[1]&INPUT_0[20]);
assign msb_1 = (INPUT_1[0]&(~INPUT_0[20])) | (comp_input1[0]&INPUT_0[20]);


assign tmp_answer[29:0] = (ans_20&{5'd30{msb_20}}) | (ans_19&{5'd30{msb_19&(~msb_20)}}) | (ans_18&{5'd30{msb_18&(~msb_19)&(~msb_20)}}) | (ans_17&{5'd30{msb_17&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_16&{5'd30{msb_16&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_15&{5'd30{msb_15&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_14&{5'd30{msb_14&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_13&{5'd30{msb_13&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_12&{5'd30{msb_12&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_11&{5'd30{msb_11&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_10&{5'd30{msb_10&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_9&{5'd30{msb_9&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_8&{5'd30{msb_8&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_7&{5'd30{msb_7&(~msb_8)&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_6&{5'd30{msb_6&(~msb_7)&(~msb_8)&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_5&{5'd30{msb_5&(~msb_6)&(~msb_7)&(~msb_8)&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_4&{5'd30{msb_4&(~msb_5)&(~msb_6)&(~msb_7)&(~msb_8)&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_3&{5'd30{msb_3&(~msb_4)&(~msb_5)&(~msb_6)&(~msb_7)&(~msb_8)&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_2&{5'd30{msb_2&(~msb_3)&(~msb_4)&(~msb_5)&(~msb_6)&(~msb_7)&(~msb_8)&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}}) | (ans_1&{5'd30{msb_1&(~msb_2)&(~msb_3)&(~msb_4)&(~msb_5)&(~msb_6)&(~msb_7)&(~msb_8)&(~msb_9)&(~msb_10)&(~msb_11)&(~msb_12)&(~msb_13)&(~msb_14)&(~msb_15)&(~msb_16)&(~msb_17)&(~msb_18)&(~msb_19)&(~msb_20)}});


assign tmp_answer[30] = 1'd0;

assign ANSWER = (tmp_answer & {5'd31{plus}}) | (((~tmp_answer)+1'd1) & {5'd31{(~plus)}});

endmodule 